
module REGISTER_FILE_NBIT64_NREG32_NADDR5 ( CLK, RST, EN, RD1, RD2, WR, DATAIN, 
        OUT1, OUT2, ADD_WR, ADD_RD1, ADD_RD2 );
  input [63:0] DATAIN;
  output [63:0] OUT1;
  output [63:0] OUT2;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input CLK, RST, EN, RD1, RD2, WR;
  wire   n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13572, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589;

  DFF_X1 \REGISTERS_reg[2][63]  ( .D(n6923), .CK(CLK), .QN(n16096) );
  DFF_X1 \REGISTERS_reg[2][62]  ( .D(n6922), .CK(CLK), .QN(n16101) );
  DFF_X1 \REGISTERS_reg[2][61]  ( .D(n6921), .CK(CLK), .QN(n16106) );
  DFF_X1 \REGISTERS_reg[2][60]  ( .D(n6920), .CK(CLK), .QN(n16111) );
  DFF_X1 \REGISTERS_reg[2][59]  ( .D(n6919), .CK(CLK), .QN(n16116) );
  DFF_X1 \REGISTERS_reg[2][58]  ( .D(n6918), .CK(CLK), .QN(n16121) );
  DFF_X1 \REGISTERS_reg[2][57]  ( .D(n6917), .CK(CLK), .QN(n16126) );
  DFF_X1 \REGISTERS_reg[2][56]  ( .D(n6916), .CK(CLK), .QN(n16131) );
  DFF_X1 \REGISTERS_reg[2][55]  ( .D(n6915), .CK(CLK), .QN(n16136) );
  DFF_X1 \REGISTERS_reg[2][54]  ( .D(n6914), .CK(CLK), .QN(n16141) );
  DFF_X1 \REGISTERS_reg[2][53]  ( .D(n6913), .CK(CLK), .QN(n16146) );
  DFF_X1 \REGISTERS_reg[2][52]  ( .D(n6912), .CK(CLK), .QN(n16151) );
  DFF_X1 \REGISTERS_reg[2][51]  ( .D(n6911), .CK(CLK), .QN(n16156) );
  DFF_X1 \REGISTERS_reg[2][50]  ( .D(n6910), .CK(CLK), .QN(n16161) );
  DFF_X1 \REGISTERS_reg[2][49]  ( .D(n6909), .CK(CLK), .QN(n16166) );
  DFF_X1 \REGISTERS_reg[2][48]  ( .D(n6908), .CK(CLK), .QN(n16171) );
  DFF_X1 \REGISTERS_reg[2][47]  ( .D(n6907), .CK(CLK), .QN(n16176) );
  DFF_X1 \REGISTERS_reg[2][46]  ( .D(n6906), .CK(CLK), .QN(n16181) );
  DFF_X1 \REGISTERS_reg[2][45]  ( .D(n6905), .CK(CLK), .QN(n16186) );
  DFF_X1 \REGISTERS_reg[2][44]  ( .D(n6904), .CK(CLK), .QN(n16191) );
  DFF_X1 \REGISTERS_reg[2][43]  ( .D(n6903), .CK(CLK), .QN(n16196) );
  DFF_X1 \REGISTERS_reg[2][42]  ( .D(n6902), .CK(CLK), .QN(n16201) );
  DFF_X1 \REGISTERS_reg[2][41]  ( .D(n6901), .CK(CLK), .QN(n16206) );
  DFF_X1 \REGISTERS_reg[2][40]  ( .D(n6900), .CK(CLK), .QN(n16211) );
  DFF_X1 \REGISTERS_reg[2][39]  ( .D(n6899), .CK(CLK), .QN(n16216) );
  DFF_X1 \REGISTERS_reg[2][38]  ( .D(n6898), .CK(CLK), .QN(n16221) );
  DFF_X1 \REGISTERS_reg[2][37]  ( .D(n6897), .CK(CLK), .QN(n16226) );
  DFF_X1 \REGISTERS_reg[2][36]  ( .D(n6896), .CK(CLK), .QN(n16231) );
  DFF_X1 \REGISTERS_reg[2][35]  ( .D(n6895), .CK(CLK), .QN(n16236) );
  DFF_X1 \REGISTERS_reg[2][34]  ( .D(n6894), .CK(CLK), .QN(n16241) );
  DFF_X1 \REGISTERS_reg[2][33]  ( .D(n6893), .CK(CLK), .QN(n16246) );
  DFF_X1 \REGISTERS_reg[2][32]  ( .D(n6892), .CK(CLK), .QN(n16251) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n6891), .CK(CLK), .QN(n16256) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n6890), .CK(CLK), .QN(n16261) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n6889), .CK(CLK), .QN(n16266) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n6888), .CK(CLK), .QN(n16271) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n6887), .CK(CLK), .QN(n16276) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n6886), .CK(CLK), .QN(n16281) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n6885), .CK(CLK), .QN(n16286) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n6884), .CK(CLK), .QN(n16291) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n6883), .CK(CLK), .QN(n16296) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n6882), .CK(CLK), .QN(n16301) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n6881), .CK(CLK), .QN(n16306) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n6880), .CK(CLK), .QN(n16311) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n6879), .CK(CLK), .QN(n16316) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n6878), .CK(CLK), .QN(n16321) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n6877), .CK(CLK), .QN(n16326) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n6876), .CK(CLK), .QN(n16331) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n6875), .CK(CLK), .QN(n16336) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n6874), .CK(CLK), .QN(n16341) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n6873), .CK(CLK), .QN(n16346) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n6872), .CK(CLK), .QN(n16351) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n6871), .CK(CLK), .QN(n16356) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n6870), .CK(CLK), .QN(n16361) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n6869), .CK(CLK), .QN(n16366) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n6868), .CK(CLK), .QN(n16371) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n6867), .CK(CLK), .QN(n16376) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n6866), .CK(CLK), .QN(n16381) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n6865), .CK(CLK), .QN(n16386) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n6864), .CK(CLK), .QN(n16391) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n6863), .CK(CLK), .QN(n16396) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n6862), .CK(CLK), .QN(n16401) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n6861), .CK(CLK), .QN(n16406) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n6860), .CK(CLK), .QN(n16411) );
  DFF_X1 \REGISTERS_reg[3][63]  ( .D(n6859), .CK(CLK), .QN(n16097) );
  DFF_X1 \REGISTERS_reg[3][62]  ( .D(n6858), .CK(CLK), .QN(n16102) );
  DFF_X1 \REGISTERS_reg[3][61]  ( .D(n6857), .CK(CLK), .QN(n16107) );
  DFF_X1 \REGISTERS_reg[3][60]  ( .D(n6856), .CK(CLK), .QN(n16112) );
  DFF_X1 \REGISTERS_reg[3][59]  ( .D(n6855), .CK(CLK), .QN(n16117) );
  DFF_X1 \REGISTERS_reg[3][58]  ( .D(n6854), .CK(CLK), .QN(n16122) );
  DFF_X1 \REGISTERS_reg[3][57]  ( .D(n6853), .CK(CLK), .QN(n16127) );
  DFF_X1 \REGISTERS_reg[3][56]  ( .D(n6852), .CK(CLK), .QN(n16132) );
  DFF_X1 \REGISTERS_reg[3][55]  ( .D(n6851), .CK(CLK), .QN(n16137) );
  DFF_X1 \REGISTERS_reg[3][54]  ( .D(n6850), .CK(CLK), .QN(n16142) );
  DFF_X1 \REGISTERS_reg[3][53]  ( .D(n6849), .CK(CLK), .QN(n16147) );
  DFF_X1 \REGISTERS_reg[3][52]  ( .D(n6848), .CK(CLK), .QN(n16152) );
  DFF_X1 \REGISTERS_reg[3][51]  ( .D(n6847), .CK(CLK), .QN(n16157) );
  DFF_X1 \REGISTERS_reg[3][50]  ( .D(n6846), .CK(CLK), .QN(n16162) );
  DFF_X1 \REGISTERS_reg[3][49]  ( .D(n6845), .CK(CLK), .QN(n16167) );
  DFF_X1 \REGISTERS_reg[3][48]  ( .D(n6844), .CK(CLK), .QN(n16172) );
  DFF_X1 \REGISTERS_reg[3][47]  ( .D(n6843), .CK(CLK), .QN(n16177) );
  DFF_X1 \REGISTERS_reg[3][46]  ( .D(n6842), .CK(CLK), .QN(n16182) );
  DFF_X1 \REGISTERS_reg[3][45]  ( .D(n6841), .CK(CLK), .QN(n16187) );
  DFF_X1 \REGISTERS_reg[3][44]  ( .D(n6840), .CK(CLK), .QN(n16192) );
  DFF_X1 \REGISTERS_reg[3][43]  ( .D(n6839), .CK(CLK), .QN(n16197) );
  DFF_X1 \REGISTERS_reg[3][42]  ( .D(n6838), .CK(CLK), .QN(n16202) );
  DFF_X1 \REGISTERS_reg[3][41]  ( .D(n6837), .CK(CLK), .QN(n16207) );
  DFF_X1 \REGISTERS_reg[3][40]  ( .D(n6836), .CK(CLK), .QN(n16212) );
  DFF_X1 \REGISTERS_reg[3][39]  ( .D(n6835), .CK(CLK), .QN(n16217) );
  DFF_X1 \REGISTERS_reg[3][38]  ( .D(n6834), .CK(CLK), .QN(n16222) );
  DFF_X1 \REGISTERS_reg[3][37]  ( .D(n6833), .CK(CLK), .QN(n16227) );
  DFF_X1 \REGISTERS_reg[3][36]  ( .D(n6832), .CK(CLK), .QN(n16232) );
  DFF_X1 \REGISTERS_reg[3][35]  ( .D(n6831), .CK(CLK), .QN(n16237) );
  DFF_X1 \REGISTERS_reg[3][34]  ( .D(n6830), .CK(CLK), .QN(n16242) );
  DFF_X1 \REGISTERS_reg[3][33]  ( .D(n6829), .CK(CLK), .QN(n16247) );
  DFF_X1 \REGISTERS_reg[3][32]  ( .D(n6828), .CK(CLK), .QN(n16252) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n6827), .CK(CLK), .QN(n16257) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n6826), .CK(CLK), .QN(n16262) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n6825), .CK(CLK), .QN(n16267) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n6824), .CK(CLK), .QN(n16272) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n6823), .CK(CLK), .QN(n16277) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n6822), .CK(CLK), .QN(n16282) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n6821), .CK(CLK), .QN(n16287) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n6820), .CK(CLK), .QN(n16292) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n6819), .CK(CLK), .QN(n16297) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n6818), .CK(CLK), .QN(n16302) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n6817), .CK(CLK), .QN(n16307) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n6816), .CK(CLK), .QN(n16312) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n6815), .CK(CLK), .QN(n16317) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n6814), .CK(CLK), .QN(n16322) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n6813), .CK(CLK), .QN(n16327) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n6812), .CK(CLK), .QN(n16332) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n6811), .CK(CLK), .QN(n16337) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n6810), .CK(CLK), .QN(n16342) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n6809), .CK(CLK), .QN(n16347) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n6808), .CK(CLK), .QN(n16352) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n6807), .CK(CLK), .QN(n16357) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n6806), .CK(CLK), .QN(n16362) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n6805), .CK(CLK), .QN(n16367) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n6804), .CK(CLK), .QN(n16372) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n6803), .CK(CLK), .QN(n16377) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n6802), .CK(CLK), .QN(n16382) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n6801), .CK(CLK), .QN(n16387) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n6800), .CK(CLK), .QN(n16392) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n6799), .CK(CLK), .QN(n16397) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n6798), .CK(CLK), .QN(n16402) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n6797), .CK(CLK), .QN(n16407) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n6796), .CK(CLK), .QN(n16412) );
  DFF_X1 \REGISTERS_reg[6][63]  ( .D(n6667), .CK(CLK), .QN(n16099) );
  DFF_X1 \REGISTERS_reg[6][62]  ( .D(n6666), .CK(CLK), .QN(n16104) );
  DFF_X1 \REGISTERS_reg[6][61]  ( .D(n6665), .CK(CLK), .QN(n16109) );
  DFF_X1 \REGISTERS_reg[6][60]  ( .D(n6664), .CK(CLK), .QN(n16114) );
  DFF_X1 \REGISTERS_reg[6][59]  ( .D(n6663), .CK(CLK), .QN(n16119) );
  DFF_X1 \REGISTERS_reg[6][58]  ( .D(n6662), .CK(CLK), .QN(n16124) );
  DFF_X1 \REGISTERS_reg[6][57]  ( .D(n6661), .CK(CLK), .QN(n16129) );
  DFF_X1 \REGISTERS_reg[6][56]  ( .D(n6660), .CK(CLK), .QN(n16134) );
  DFF_X1 \REGISTERS_reg[6][55]  ( .D(n6659), .CK(CLK), .QN(n16139) );
  DFF_X1 \REGISTERS_reg[6][54]  ( .D(n6658), .CK(CLK), .QN(n16144) );
  DFF_X1 \REGISTERS_reg[6][53]  ( .D(n6657), .CK(CLK), .QN(n16149) );
  DFF_X1 \REGISTERS_reg[6][52]  ( .D(n6656), .CK(CLK), .QN(n16154) );
  DFF_X1 \REGISTERS_reg[6][51]  ( .D(n6655), .CK(CLK), .QN(n16159) );
  DFF_X1 \REGISTERS_reg[6][50]  ( .D(n6654), .CK(CLK), .QN(n16164) );
  DFF_X1 \REGISTERS_reg[6][49]  ( .D(n6653), .CK(CLK), .QN(n16169) );
  DFF_X1 \REGISTERS_reg[6][48]  ( .D(n6652), .CK(CLK), .QN(n16174) );
  DFF_X1 \REGISTERS_reg[6][47]  ( .D(n6651), .CK(CLK), .QN(n16179) );
  DFF_X1 \REGISTERS_reg[6][46]  ( .D(n6650), .CK(CLK), .QN(n16184) );
  DFF_X1 \REGISTERS_reg[6][45]  ( .D(n6649), .CK(CLK), .QN(n16189) );
  DFF_X1 \REGISTERS_reg[6][44]  ( .D(n6648), .CK(CLK), .QN(n16194) );
  DFF_X1 \REGISTERS_reg[6][43]  ( .D(n6647), .CK(CLK), .QN(n16199) );
  DFF_X1 \REGISTERS_reg[6][42]  ( .D(n6646), .CK(CLK), .QN(n16204) );
  DFF_X1 \REGISTERS_reg[6][41]  ( .D(n6645), .CK(CLK), .QN(n16209) );
  DFF_X1 \REGISTERS_reg[6][40]  ( .D(n6644), .CK(CLK), .QN(n16214) );
  DFF_X1 \REGISTERS_reg[6][39]  ( .D(n6643), .CK(CLK), .QN(n16219) );
  DFF_X1 \REGISTERS_reg[6][38]  ( .D(n6642), .CK(CLK), .QN(n16224) );
  DFF_X1 \REGISTERS_reg[6][37]  ( .D(n6641), .CK(CLK), .QN(n16229) );
  DFF_X1 \REGISTERS_reg[6][36]  ( .D(n6640), .CK(CLK), .QN(n16234) );
  DFF_X1 \REGISTERS_reg[6][35]  ( .D(n6639), .CK(CLK), .QN(n16239) );
  DFF_X1 \REGISTERS_reg[6][34]  ( .D(n6638), .CK(CLK), .QN(n16244) );
  DFF_X1 \REGISTERS_reg[6][33]  ( .D(n6637), .CK(CLK), .QN(n16249) );
  DFF_X1 \REGISTERS_reg[6][32]  ( .D(n6636), .CK(CLK), .QN(n16254) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n6635), .CK(CLK), .QN(n16259) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n6634), .CK(CLK), .QN(n16264) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n6633), .CK(CLK), .QN(n16269) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n6632), .CK(CLK), .QN(n16274) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n6631), .CK(CLK), .QN(n16279) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n6630), .CK(CLK), .QN(n16284) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n6629), .CK(CLK), .QN(n16289) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n6628), .CK(CLK), .QN(n16294) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n6627), .CK(CLK), .QN(n16299) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n6626), .CK(CLK), .QN(n16304) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n6625), .CK(CLK), .QN(n16309) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n6624), .CK(CLK), .QN(n16314) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n6623), .CK(CLK), .QN(n16319) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n6622), .CK(CLK), .QN(n16324) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n6621), .CK(CLK), .QN(n16329) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n6620), .CK(CLK), .QN(n16334) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n6619), .CK(CLK), .QN(n16339) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n6618), .CK(CLK), .QN(n16344) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n6617), .CK(CLK), .QN(n16349) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n6616), .CK(CLK), .QN(n16354) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n6615), .CK(CLK), .QN(n16359) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n6614), .CK(CLK), .QN(n16364) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n6613), .CK(CLK), .QN(n16369) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n6612), .CK(CLK), .QN(n16374) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n6611), .CK(CLK), .QN(n16379) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n6610), .CK(CLK), .QN(n16384) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n6609), .CK(CLK), .QN(n16389) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n6608), .CK(CLK), .QN(n16394) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n6607), .CK(CLK), .QN(n16399) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n6606), .CK(CLK), .QN(n16404) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n6605), .CK(CLK), .QN(n16409) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n6604), .CK(CLK), .QN(n16414) );
  DFF_X1 \REGISTERS_reg[7][63]  ( .D(n6603), .CK(CLK), .QN(n16098) );
  DFF_X1 \REGISTERS_reg[7][62]  ( .D(n6602), .CK(CLK), .QN(n16103) );
  DFF_X1 \REGISTERS_reg[7][61]  ( .D(n6601), .CK(CLK), .QN(n16108) );
  DFF_X1 \REGISTERS_reg[7][60]  ( .D(n6600), .CK(CLK), .QN(n16113) );
  DFF_X1 \REGISTERS_reg[7][59]  ( .D(n6599), .CK(CLK), .QN(n16118) );
  DFF_X1 \REGISTERS_reg[7][58]  ( .D(n6598), .CK(CLK), .QN(n16123) );
  DFF_X1 \REGISTERS_reg[7][57]  ( .D(n6597), .CK(CLK), .QN(n16128) );
  DFF_X1 \REGISTERS_reg[7][56]  ( .D(n6596), .CK(CLK), .QN(n16133) );
  DFF_X1 \REGISTERS_reg[7][55]  ( .D(n6595), .CK(CLK), .QN(n16138) );
  DFF_X1 \REGISTERS_reg[7][54]  ( .D(n6594), .CK(CLK), .QN(n16143) );
  DFF_X1 \REGISTERS_reg[7][53]  ( .D(n6593), .CK(CLK), .QN(n16148) );
  DFF_X1 \REGISTERS_reg[7][52]  ( .D(n6592), .CK(CLK), .QN(n16153) );
  DFF_X1 \REGISTERS_reg[7][51]  ( .D(n6591), .CK(CLK), .QN(n16158) );
  DFF_X1 \REGISTERS_reg[7][50]  ( .D(n6590), .CK(CLK), .QN(n16163) );
  DFF_X1 \REGISTERS_reg[7][49]  ( .D(n6589), .CK(CLK), .QN(n16168) );
  DFF_X1 \REGISTERS_reg[7][48]  ( .D(n6588), .CK(CLK), .QN(n16173) );
  DFF_X1 \REGISTERS_reg[7][47]  ( .D(n6587), .CK(CLK), .QN(n16178) );
  DFF_X1 \REGISTERS_reg[7][46]  ( .D(n6586), .CK(CLK), .QN(n16183) );
  DFF_X1 \REGISTERS_reg[7][45]  ( .D(n6585), .CK(CLK), .QN(n16188) );
  DFF_X1 \REGISTERS_reg[7][44]  ( .D(n6584), .CK(CLK), .QN(n16193) );
  DFF_X1 \REGISTERS_reg[7][43]  ( .D(n6583), .CK(CLK), .QN(n16198) );
  DFF_X1 \REGISTERS_reg[7][42]  ( .D(n6582), .CK(CLK), .QN(n16203) );
  DFF_X1 \REGISTERS_reg[7][41]  ( .D(n6581), .CK(CLK), .QN(n16208) );
  DFF_X1 \REGISTERS_reg[7][40]  ( .D(n6580), .CK(CLK), .QN(n16213) );
  DFF_X1 \REGISTERS_reg[7][39]  ( .D(n6579), .CK(CLK), .QN(n16218) );
  DFF_X1 \REGISTERS_reg[7][38]  ( .D(n6578), .CK(CLK), .QN(n16223) );
  DFF_X1 \REGISTERS_reg[7][37]  ( .D(n6577), .CK(CLK), .QN(n16228) );
  DFF_X1 \REGISTERS_reg[7][36]  ( .D(n6576), .CK(CLK), .QN(n16233) );
  DFF_X1 \REGISTERS_reg[7][35]  ( .D(n6575), .CK(CLK), .QN(n16238) );
  DFF_X1 \REGISTERS_reg[7][34]  ( .D(n6574), .CK(CLK), .QN(n16243) );
  DFF_X1 \REGISTERS_reg[7][33]  ( .D(n6573), .CK(CLK), .QN(n16248) );
  DFF_X1 \REGISTERS_reg[7][32]  ( .D(n6572), .CK(CLK), .QN(n16253) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n6571), .CK(CLK), .QN(n16258) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n6570), .CK(CLK), .QN(n16263) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n6569), .CK(CLK), .QN(n16268) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n6568), .CK(CLK), .QN(n16273) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n6567), .CK(CLK), .QN(n16278) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n6566), .CK(CLK), .QN(n16283) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n6565), .CK(CLK), .QN(n16288) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n6564), .CK(CLK), .QN(n16293) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n6563), .CK(CLK), .QN(n16298) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n6562), .CK(CLK), .QN(n16303) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n6561), .CK(CLK), .QN(n16308) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n6560), .CK(CLK), .QN(n16313) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n6559), .CK(CLK), .QN(n16318) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n6558), .CK(CLK), .QN(n16323) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n6557), .CK(CLK), .QN(n16328) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n6556), .CK(CLK), .QN(n16333) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n6555), .CK(CLK), .QN(n16338) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n6554), .CK(CLK), .QN(n16343) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n6553), .CK(CLK), .QN(n16348) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n6552), .CK(CLK), .QN(n16353) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n6551), .CK(CLK), .QN(n16358) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n6550), .CK(CLK), .QN(n16363) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n6549), .CK(CLK), .QN(n16368) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n6548), .CK(CLK), .QN(n16373) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n6547), .CK(CLK), .QN(n16378) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n6546), .CK(CLK), .QN(n16383) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n6545), .CK(CLK), .QN(n16388) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n6544), .CK(CLK), .QN(n16393) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n6543), .CK(CLK), .QN(n16398) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n6542), .CK(CLK), .QN(n16403) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n6541), .CK(CLK), .QN(n16408) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n6540), .CK(CLK), .QN(n16413) );
  DFF_X1 \REGISTERS_reg[13][63]  ( .D(n6219), .CK(CLK), .QN(n837) );
  DFF_X1 \REGISTERS_reg[13][62]  ( .D(n6218), .CK(CLK), .QN(n838) );
  DFF_X1 \REGISTERS_reg[13][61]  ( .D(n6217), .CK(CLK), .QN(n839) );
  DFF_X1 \REGISTERS_reg[13][60]  ( .D(n6216), .CK(CLK), .QN(n840) );
  DFF_X1 \REGISTERS_reg[13][59]  ( .D(n6215), .CK(CLK), .QN(n841) );
  DFF_X1 \REGISTERS_reg[13][58]  ( .D(n6214), .CK(CLK), .QN(n842) );
  DFF_X1 \REGISTERS_reg[13][57]  ( .D(n6213), .CK(CLK), .QN(n843) );
  DFF_X1 \REGISTERS_reg[13][56]  ( .D(n6212), .CK(CLK), .QN(n844) );
  DFF_X1 \REGISTERS_reg[13][55]  ( .D(n6211), .CK(CLK), .QN(n845) );
  DFF_X1 \REGISTERS_reg[13][54]  ( .D(n6210), .CK(CLK), .QN(n846) );
  DFF_X1 \REGISTERS_reg[13][53]  ( .D(n6209), .CK(CLK), .QN(n847) );
  DFF_X1 \REGISTERS_reg[13][52]  ( .D(n6208), .CK(CLK), .QN(n848) );
  DFF_X1 \REGISTERS_reg[13][51]  ( .D(n6207), .CK(CLK), .QN(n849) );
  DFF_X1 \REGISTERS_reg[13][50]  ( .D(n6206), .CK(CLK), .QN(n850) );
  DFF_X1 \REGISTERS_reg[13][49]  ( .D(n6205), .CK(CLK), .QN(n851) );
  DFF_X1 \REGISTERS_reg[13][48]  ( .D(n6204), .CK(CLK), .QN(n852) );
  DFF_X1 \REGISTERS_reg[13][47]  ( .D(n6203), .CK(CLK), .QN(n853) );
  DFF_X1 \REGISTERS_reg[13][46]  ( .D(n6202), .CK(CLK), .QN(n854) );
  DFF_X1 \REGISTERS_reg[13][45]  ( .D(n6201), .CK(CLK), .QN(n855) );
  DFF_X1 \REGISTERS_reg[13][44]  ( .D(n6200), .CK(CLK), .QN(n856) );
  DFF_X1 \REGISTERS_reg[13][43]  ( .D(n6199), .CK(CLK), .QN(n857) );
  DFF_X1 \REGISTERS_reg[13][42]  ( .D(n6198), .CK(CLK), .QN(n858) );
  DFF_X1 \REGISTERS_reg[13][41]  ( .D(n6197), .CK(CLK), .QN(n859) );
  DFF_X1 \REGISTERS_reg[13][40]  ( .D(n6196), .CK(CLK), .QN(n860) );
  DFF_X1 \REGISTERS_reg[13][39]  ( .D(n6195), .CK(CLK), .QN(n861) );
  DFF_X1 \REGISTERS_reg[13][38]  ( .D(n6194), .CK(CLK), .QN(n862) );
  DFF_X1 \REGISTERS_reg[13][37]  ( .D(n6193), .CK(CLK), .QN(n863) );
  DFF_X1 \REGISTERS_reg[13][36]  ( .D(n6192), .CK(CLK), .QN(n864) );
  DFF_X1 \REGISTERS_reg[13][35]  ( .D(n6191), .CK(CLK), .QN(n865) );
  DFF_X1 \REGISTERS_reg[13][34]  ( .D(n6190), .CK(CLK), .QN(n866) );
  DFF_X1 \REGISTERS_reg[13][33]  ( .D(n6189), .CK(CLK), .QN(n867) );
  DFF_X1 \REGISTERS_reg[13][32]  ( .D(n6188), .CK(CLK), .QN(n868) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n6187), .CK(CLK), .QN(n869) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n6186), .CK(CLK), .QN(n870) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n6185), .CK(CLK), .QN(n871) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n6184), .CK(CLK), .QN(n872) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n6183), .CK(CLK), .QN(n873) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n6182), .CK(CLK), .QN(n874) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n6181), .CK(CLK), .QN(n875) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n6180), .CK(CLK), .QN(n876) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n6179), .CK(CLK), .QN(n877) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n6178), .CK(CLK), .QN(n878) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n6177), .CK(CLK), .QN(n879) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n6176), .CK(CLK), .QN(n880) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n6175), .CK(CLK), .QN(n881) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n6174), .CK(CLK), .QN(n882) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n6173), .CK(CLK), .QN(n883) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n6172), .CK(CLK), .QN(n884) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n6171), .CK(CLK), .QN(n885) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n6170), .CK(CLK), .QN(n886) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n6169), .CK(CLK), .QN(n887) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n6168), .CK(CLK), .QN(n888) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n6167), .CK(CLK), .QN(n889) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n6166), .CK(CLK), .QN(n890) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n6165), .CK(CLK), .QN(n891) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n6164), .CK(CLK), .QN(n892) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n6163), .CK(CLK), .QN(n893) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n6162), .CK(CLK), .QN(n894) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n6161), .CK(CLK), .QN(n895) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n6160), .CK(CLK), .QN(n896) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n6159), .CK(CLK), .QN(n897) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n6158), .CK(CLK), .QN(n898) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n6157), .CK(CLK), .QN(n899) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n6156), .CK(CLK), .QN(n900) );
  DFF_X1 \REGISTERS_reg[14][63]  ( .D(n6155), .CK(CLK), .QN(n901) );
  DFF_X1 \REGISTERS_reg[14][62]  ( .D(n6154), .CK(CLK), .QN(n902) );
  DFF_X1 \REGISTERS_reg[14][61]  ( .D(n6153), .CK(CLK), .QN(n903) );
  DFF_X1 \REGISTERS_reg[14][60]  ( .D(n6152), .CK(CLK), .QN(n904) );
  DFF_X1 \REGISTERS_reg[14][59]  ( .D(n6151), .CK(CLK), .QN(n905) );
  DFF_X1 \REGISTERS_reg[14][58]  ( .D(n6150), .CK(CLK), .QN(n906) );
  DFF_X1 \REGISTERS_reg[14][57]  ( .D(n6149), .CK(CLK), .QN(n907) );
  DFF_X1 \REGISTERS_reg[14][56]  ( .D(n6148), .CK(CLK), .QN(n908) );
  DFF_X1 \REGISTERS_reg[14][55]  ( .D(n6147), .CK(CLK), .QN(n909) );
  DFF_X1 \REGISTERS_reg[14][54]  ( .D(n6146), .CK(CLK), .QN(n910) );
  DFF_X1 \REGISTERS_reg[14][53]  ( .D(n6145), .CK(CLK), .QN(n911) );
  DFF_X1 \REGISTERS_reg[14][52]  ( .D(n6144), .CK(CLK), .QN(n912) );
  DFF_X1 \REGISTERS_reg[14][51]  ( .D(n6143), .CK(CLK), .QN(n913) );
  DFF_X1 \REGISTERS_reg[14][50]  ( .D(n6142), .CK(CLK), .QN(n914) );
  DFF_X1 \REGISTERS_reg[14][49]  ( .D(n6141), .CK(CLK), .QN(n915) );
  DFF_X1 \REGISTERS_reg[14][48]  ( .D(n6140), .CK(CLK), .QN(n916) );
  DFF_X1 \REGISTERS_reg[14][47]  ( .D(n6139), .CK(CLK), .QN(n917) );
  DFF_X1 \REGISTERS_reg[14][46]  ( .D(n6138), .CK(CLK), .QN(n918) );
  DFF_X1 \REGISTERS_reg[14][45]  ( .D(n6137), .CK(CLK), .QN(n919) );
  DFF_X1 \REGISTERS_reg[14][44]  ( .D(n6136), .CK(CLK), .QN(n920) );
  DFF_X1 \REGISTERS_reg[14][43]  ( .D(n6135), .CK(CLK), .QN(n921) );
  DFF_X1 \REGISTERS_reg[14][42]  ( .D(n6134), .CK(CLK), .QN(n922) );
  DFF_X1 \REGISTERS_reg[14][41]  ( .D(n6133), .CK(CLK), .QN(n923) );
  DFF_X1 \REGISTERS_reg[14][40]  ( .D(n6132), .CK(CLK), .QN(n924) );
  DFF_X1 \REGISTERS_reg[14][39]  ( .D(n6131), .CK(CLK), .QN(n925) );
  DFF_X1 \REGISTERS_reg[14][38]  ( .D(n6130), .CK(CLK), .QN(n926) );
  DFF_X1 \REGISTERS_reg[14][37]  ( .D(n6129), .CK(CLK), .QN(n927) );
  DFF_X1 \REGISTERS_reg[14][36]  ( .D(n6128), .CK(CLK), .QN(n928) );
  DFF_X1 \REGISTERS_reg[14][35]  ( .D(n6127), .CK(CLK), .QN(n929) );
  DFF_X1 \REGISTERS_reg[14][34]  ( .D(n6126), .CK(CLK), .QN(n930) );
  DFF_X1 \REGISTERS_reg[14][33]  ( .D(n6125), .CK(CLK), .QN(n931) );
  DFF_X1 \REGISTERS_reg[14][32]  ( .D(n6124), .CK(CLK), .QN(n932) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n6123), .CK(CLK), .QN(n933) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n6122), .CK(CLK), .QN(n934) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n6121), .CK(CLK), .QN(n935) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n6120), .CK(CLK), .QN(n936) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n6119), .CK(CLK), .QN(n937) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n6118), .CK(CLK), .QN(n938) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n6117), .CK(CLK), .QN(n939) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n6116), .CK(CLK), .QN(n940) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n6115), .CK(CLK), .QN(n941) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n6114), .CK(CLK), .QN(n942) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n6113), .CK(CLK), .QN(n943) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n6112), .CK(CLK), .QN(n944) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n6111), .CK(CLK), .QN(n945) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n6110), .CK(CLK), .QN(n946) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n6109), .CK(CLK), .QN(n947) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n6108), .CK(CLK), .QN(n948) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n6107), .CK(CLK), .QN(n949) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n6106), .CK(CLK), .QN(n950) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n6105), .CK(CLK), .QN(n951) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n6104), .CK(CLK), .QN(n952) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n6103), .CK(CLK), .QN(n953) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n6102), .CK(CLK), .QN(n954) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n6101), .CK(CLK), .QN(n955) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n6100), .CK(CLK), .QN(n956) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n6099), .CK(CLK), .QN(n957) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n6098), .CK(CLK), .QN(n958) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n6097), .CK(CLK), .QN(n959) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n6096), .CK(CLK), .QN(n960) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n6095), .CK(CLK), .QN(n961) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n6094), .CK(CLK), .QN(n962) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n6093), .CK(CLK), .QN(n963) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n6092), .CK(CLK), .QN(n964) );
  DFF_X1 \REGISTERS_reg[15][63]  ( .D(n6091), .CK(CLK), .QN(n965) );
  DFF_X1 \REGISTERS_reg[15][62]  ( .D(n6090), .CK(CLK), .QN(n966) );
  DFF_X1 \REGISTERS_reg[15][61]  ( .D(n6089), .CK(CLK), .QN(n967) );
  DFF_X1 \REGISTERS_reg[15][60]  ( .D(n6088), .CK(CLK), .QN(n968) );
  DFF_X1 \REGISTERS_reg[15][59]  ( .D(n6087), .CK(CLK), .QN(n969) );
  DFF_X1 \REGISTERS_reg[15][58]  ( .D(n6086), .CK(CLK), .QN(n970) );
  DFF_X1 \REGISTERS_reg[15][57]  ( .D(n6085), .CK(CLK), .QN(n971) );
  DFF_X1 \REGISTERS_reg[15][56]  ( .D(n6084), .CK(CLK), .QN(n972) );
  DFF_X1 \REGISTERS_reg[15][55]  ( .D(n6083), .CK(CLK), .QN(n973) );
  DFF_X1 \REGISTERS_reg[15][54]  ( .D(n6082), .CK(CLK), .QN(n974) );
  DFF_X1 \REGISTERS_reg[15][53]  ( .D(n6081), .CK(CLK), .QN(n975) );
  DFF_X1 \REGISTERS_reg[15][52]  ( .D(n6080), .CK(CLK), .QN(n976) );
  DFF_X1 \REGISTERS_reg[15][51]  ( .D(n6079), .CK(CLK), .QN(n977) );
  DFF_X1 \REGISTERS_reg[15][50]  ( .D(n6078), .CK(CLK), .QN(n978) );
  DFF_X1 \REGISTERS_reg[15][49]  ( .D(n6077), .CK(CLK), .QN(n979) );
  DFF_X1 \REGISTERS_reg[15][48]  ( .D(n6076), .CK(CLK), .QN(n980) );
  DFF_X1 \REGISTERS_reg[15][47]  ( .D(n6075), .CK(CLK), .QN(n981) );
  DFF_X1 \REGISTERS_reg[15][46]  ( .D(n6074), .CK(CLK), .QN(n982) );
  DFF_X1 \REGISTERS_reg[15][45]  ( .D(n6073), .CK(CLK), .QN(n983) );
  DFF_X1 \REGISTERS_reg[15][44]  ( .D(n6072), .CK(CLK), .QN(n984) );
  DFF_X1 \REGISTERS_reg[15][43]  ( .D(n6071), .CK(CLK), .QN(n985) );
  DFF_X1 \REGISTERS_reg[15][42]  ( .D(n6070), .CK(CLK), .QN(n986) );
  DFF_X1 \REGISTERS_reg[15][41]  ( .D(n6069), .CK(CLK), .QN(n987) );
  DFF_X1 \REGISTERS_reg[15][40]  ( .D(n6068), .CK(CLK), .QN(n988) );
  DFF_X1 \REGISTERS_reg[15][39]  ( .D(n6067), .CK(CLK), .QN(n989) );
  DFF_X1 \REGISTERS_reg[15][38]  ( .D(n6066), .CK(CLK), .QN(n990) );
  DFF_X1 \REGISTERS_reg[15][37]  ( .D(n6065), .CK(CLK), .QN(n991) );
  DFF_X1 \REGISTERS_reg[15][36]  ( .D(n6064), .CK(CLK), .QN(n992) );
  DFF_X1 \REGISTERS_reg[15][35]  ( .D(n6063), .CK(CLK), .QN(n993) );
  DFF_X1 \REGISTERS_reg[15][34]  ( .D(n6062), .CK(CLK), .QN(n994) );
  DFF_X1 \REGISTERS_reg[15][33]  ( .D(n6061), .CK(CLK), .QN(n995) );
  DFF_X1 \REGISTERS_reg[15][32]  ( .D(n6060), .CK(CLK), .QN(n996) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n6059), .CK(CLK), .QN(n997) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n6058), .CK(CLK), .QN(n998) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n6057), .CK(CLK), .QN(n999) );
  DFF_X1 \REGISTERS_reg[18][63]  ( .D(n5899), .CK(CLK), .QN(n7610) );
  DFF_X1 \REGISTERS_reg[18][62]  ( .D(n5898), .CK(CLK), .QN(n7612) );
  DFF_X1 \REGISTERS_reg[18][61]  ( .D(n5897), .CK(CLK), .QN(n7614) );
  DFF_X1 \REGISTERS_reg[18][60]  ( .D(n5896), .CK(CLK), .QN(n7616) );
  DFF_X1 \REGISTERS_reg[18][59]  ( .D(n5895), .CK(CLK), .QN(n7618) );
  DFF_X1 \REGISTERS_reg[18][58]  ( .D(n5894), .CK(CLK), .QN(n7620) );
  DFF_X1 \REGISTERS_reg[18][57]  ( .D(n5893), .CK(CLK), .QN(n7622) );
  DFF_X1 \REGISTERS_reg[18][56]  ( .D(n5892), .CK(CLK), .QN(n7624) );
  DFF_X1 \REGISTERS_reg[18][55]  ( .D(n5891), .CK(CLK), .QN(n7626) );
  DFF_X1 \REGISTERS_reg[18][54]  ( .D(n5890), .CK(CLK), .QN(n7628) );
  DFF_X1 \REGISTERS_reg[18][53]  ( .D(n5889), .CK(CLK), .QN(n7630) );
  DFF_X1 \REGISTERS_reg[18][52]  ( .D(n5888), .CK(CLK), .QN(n7632) );
  DFF_X1 \REGISTERS_reg[18][51]  ( .D(n5887), .CK(CLK), .QN(n7634) );
  DFF_X1 \REGISTERS_reg[18][50]  ( .D(n5886), .CK(CLK), .QN(n7636) );
  DFF_X1 \REGISTERS_reg[18][49]  ( .D(n5885), .CK(CLK), .QN(n7638) );
  DFF_X1 \REGISTERS_reg[18][48]  ( .D(n5884), .CK(CLK), .QN(n7640) );
  DFF_X1 \REGISTERS_reg[18][47]  ( .D(n5883), .CK(CLK), .QN(n7642) );
  DFF_X1 \REGISTERS_reg[18][46]  ( .D(n5882), .CK(CLK), .QN(n7644) );
  DFF_X1 \REGISTERS_reg[18][45]  ( .D(n5881), .CK(CLK), .QN(n7646) );
  DFF_X1 \REGISTERS_reg[18][44]  ( .D(n5880), .CK(CLK), .QN(n7648) );
  DFF_X1 \REGISTERS_reg[18][43]  ( .D(n5879), .CK(CLK), .QN(n7650) );
  DFF_X1 \REGISTERS_reg[18][42]  ( .D(n5878), .CK(CLK), .QN(n7652) );
  DFF_X1 \REGISTERS_reg[18][41]  ( .D(n5877), .CK(CLK), .QN(n7654) );
  DFF_X1 \REGISTERS_reg[18][40]  ( .D(n5876), .CK(CLK), .QN(n7656) );
  DFF_X1 \REGISTERS_reg[18][39]  ( .D(n5875), .CK(CLK), .QN(n7658) );
  DFF_X1 \REGISTERS_reg[18][38]  ( .D(n5874), .CK(CLK), .QN(n7660) );
  DFF_X1 \REGISTERS_reg[18][37]  ( .D(n5873), .CK(CLK), .QN(n7662) );
  DFF_X1 \REGISTERS_reg[18][36]  ( .D(n5872), .CK(CLK), .QN(n7664) );
  DFF_X1 \REGISTERS_reg[18][35]  ( .D(n5871), .CK(CLK), .QN(n7666) );
  DFF_X1 \REGISTERS_reg[18][34]  ( .D(n5870), .CK(CLK), .QN(n7668) );
  DFF_X1 \REGISTERS_reg[18][33]  ( .D(n5869), .CK(CLK), .QN(n7670) );
  DFF_X1 \REGISTERS_reg[18][32]  ( .D(n5868), .CK(CLK), .QN(n7672) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n5867), .CK(CLK), .QN(n7674) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n5866), .CK(CLK), .QN(n7676) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n5865), .CK(CLK), .QN(n7678) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n5864), .CK(CLK), .QN(n7680) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n5863), .CK(CLK), .QN(n7682) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n5862), .CK(CLK), .QN(n7684) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n5861), .CK(CLK), .QN(n7686) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n5860), .CK(CLK), .QN(n7688) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n5859), .CK(CLK), .QN(n7690) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n5858), .CK(CLK), .QN(n7692) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n5857), .CK(CLK), .QN(n7694) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n5856), .CK(CLK), .QN(n7696) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n5855), .CK(CLK), .QN(n7698) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n5854), .CK(CLK), .QN(n7700) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n5853), .CK(CLK), .QN(n7702) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n5852), .CK(CLK), .QN(n7704) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n5851), .CK(CLK), .QN(n7706) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n5850), .CK(CLK), .QN(n7708) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n5849), .CK(CLK), .QN(n7710) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n5848), .CK(CLK), .QN(n7712) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n5847), .CK(CLK), .QN(n7714) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n5846), .CK(CLK), .QN(n7716) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n5845), .CK(CLK), .QN(n7718) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n5844), .CK(CLK), .QN(n7720) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n5843), .CK(CLK), .QN(n7722) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n5842), .CK(CLK), .QN(n7724) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n5841), .CK(CLK), .QN(n7726) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n5840), .CK(CLK), .QN(n7728) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n5839), .CK(CLK), .QN(n7730) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n5838), .CK(CLK), .QN(n7732) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n5837), .CK(CLK), .QN(n7734) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n5836), .CK(CLK), .QN(n7736) );
  DFF_X1 \REGISTERS_reg[19][63]  ( .D(n5835), .CK(CLK), .QN(n7738) );
  DFF_X1 \REGISTERS_reg[19][62]  ( .D(n5834), .CK(CLK), .QN(n7740) );
  DFF_X1 \REGISTERS_reg[19][61]  ( .D(n5833), .CK(CLK), .QN(n7742) );
  DFF_X1 \REGISTERS_reg[19][60]  ( .D(n5832), .CK(CLK), .QN(n7744) );
  DFF_X1 \REGISTERS_reg[19][59]  ( .D(n5831), .CK(CLK), .QN(n7746) );
  DFF_X1 \REGISTERS_reg[19][58]  ( .D(n5830), .CK(CLK), .QN(n7748) );
  DFF_X1 \REGISTERS_reg[19][57]  ( .D(n5829), .CK(CLK), .QN(n7750) );
  DFF_X1 \REGISTERS_reg[19][56]  ( .D(n5828), .CK(CLK), .QN(n7752) );
  DFF_X1 \REGISTERS_reg[19][55]  ( .D(n5827), .CK(CLK), .QN(n7754) );
  DFF_X1 \REGISTERS_reg[19][54]  ( .D(n5826), .CK(CLK), .QN(n7756) );
  DFF_X1 \REGISTERS_reg[19][53]  ( .D(n5825), .CK(CLK), .QN(n7758) );
  DFF_X1 \REGISTERS_reg[19][52]  ( .D(n5824), .CK(CLK), .QN(n7760) );
  DFF_X1 \REGISTERS_reg[19][51]  ( .D(n5823), .CK(CLK), .QN(n7762) );
  DFF_X1 \REGISTERS_reg[19][50]  ( .D(n5822), .CK(CLK), .QN(n7764) );
  DFF_X1 \REGISTERS_reg[19][49]  ( .D(n5821), .CK(CLK), .QN(n7766) );
  DFF_X1 \REGISTERS_reg[19][48]  ( .D(n5820), .CK(CLK), .QN(n7768) );
  DFF_X1 \REGISTERS_reg[19][47]  ( .D(n5819), .CK(CLK), .QN(n7770) );
  DFF_X1 \REGISTERS_reg[19][46]  ( .D(n5818), .CK(CLK), .QN(n7772) );
  DFF_X1 \REGISTERS_reg[19][45]  ( .D(n5817), .CK(CLK), .QN(n7774) );
  DFF_X1 \REGISTERS_reg[19][44]  ( .D(n5816), .CK(CLK), .QN(n7776) );
  DFF_X1 \REGISTERS_reg[19][43]  ( .D(n5815), .CK(CLK), .QN(n7778) );
  DFF_X1 \REGISTERS_reg[19][42]  ( .D(n5814), .CK(CLK), .QN(n7780) );
  DFF_X1 \REGISTERS_reg[19][41]  ( .D(n5813), .CK(CLK), .QN(n7782) );
  DFF_X1 \REGISTERS_reg[19][40]  ( .D(n5812), .CK(CLK), .QN(n7784) );
  DFF_X1 \REGISTERS_reg[19][39]  ( .D(n5811), .CK(CLK), .QN(n7786) );
  DFF_X1 \REGISTERS_reg[19][38]  ( .D(n5810), .CK(CLK), .QN(n7788) );
  DFF_X1 \REGISTERS_reg[19][37]  ( .D(n5809), .CK(CLK), .QN(n7790) );
  DFF_X1 \REGISTERS_reg[19][36]  ( .D(n5808), .CK(CLK), .QN(n7792) );
  DFF_X1 \REGISTERS_reg[19][35]  ( .D(n5807), .CK(CLK), .QN(n7794) );
  DFF_X1 \REGISTERS_reg[19][34]  ( .D(n5806), .CK(CLK), .QN(n7796) );
  DFF_X1 \REGISTERS_reg[19][33]  ( .D(n5805), .CK(CLK), .QN(n7798) );
  DFF_X1 \REGISTERS_reg[19][32]  ( .D(n5804), .CK(CLK), .QN(n7800) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n5803), .CK(CLK), .QN(n7802) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n5802), .CK(CLK), .QN(n7804) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n5801), .CK(CLK), .QN(n7806) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n5800), .CK(CLK), .QN(n7808) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n5799), .CK(CLK), .QN(n7810) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n5798), .CK(CLK), .QN(n7812) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n5797), .CK(CLK), .QN(n7814) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n5796), .CK(CLK), .QN(n7816) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n5795), .CK(CLK), .QN(n7818) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n5794), .CK(CLK), .QN(n7820) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n5793), .CK(CLK), .QN(n7822) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n5792), .CK(CLK), .QN(n7824) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n5791), .CK(CLK), .QN(n7826) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n5790), .CK(CLK), .QN(n7828) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n5789), .CK(CLK), .QN(n7830) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n5788), .CK(CLK), .QN(n7832) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n5787), .CK(CLK), .QN(n7834) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n5786), .CK(CLK), .QN(n7836) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n5785), .CK(CLK), .QN(n7838) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n5784), .CK(CLK), .QN(n7840) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n5783), .CK(CLK), .QN(n7842) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n5782), .CK(CLK), .QN(n7844) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n5781), .CK(CLK), .QN(n7846) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n5780), .CK(CLK), .QN(n7848) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n5779), .CK(CLK), .QN(n7850) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n5778), .CK(CLK), .QN(n7852) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n5777), .CK(CLK), .QN(n7854) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n5776), .CK(CLK), .QN(n7856) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n5775), .CK(CLK), .QN(n7858) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n5774), .CK(CLK), .QN(n7860) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n5773), .CK(CLK), .QN(n7862) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n5772), .CK(CLK), .QN(n7864) );
  DFF_X1 \REGISTERS_reg[23][63]  ( .D(n5579), .CK(CLK), .QN(n7866) );
  DFF_X1 \REGISTERS_reg[23][62]  ( .D(n5578), .CK(CLK), .QN(n7869) );
  DFF_X1 \REGISTERS_reg[23][61]  ( .D(n5577), .CK(CLK), .QN(n7872) );
  DFF_X1 \REGISTERS_reg[23][60]  ( .D(n5576), .CK(CLK), .QN(n7875) );
  DFF_X1 \REGISTERS_reg[23][59]  ( .D(n5575), .CK(CLK), .QN(n7878) );
  DFF_X1 \REGISTERS_reg[23][58]  ( .D(n5574), .CK(CLK), .QN(n7881) );
  DFF_X1 \REGISTERS_reg[23][57]  ( .D(n5573), .CK(CLK), .QN(n7884) );
  DFF_X1 \REGISTERS_reg[23][56]  ( .D(n5572), .CK(CLK), .QN(n7887) );
  DFF_X1 \REGISTERS_reg[23][55]  ( .D(n5571), .CK(CLK), .QN(n7890) );
  DFF_X1 \REGISTERS_reg[23][54]  ( .D(n5570), .CK(CLK), .QN(n7893) );
  DFF_X1 \REGISTERS_reg[23][53]  ( .D(n5569), .CK(CLK), .QN(n7896) );
  DFF_X1 \REGISTERS_reg[23][52]  ( .D(n5568), .CK(CLK), .QN(n7899) );
  DFF_X1 \REGISTERS_reg[23][51]  ( .D(n5567), .CK(CLK), .QN(n7902) );
  DFF_X1 \REGISTERS_reg[23][50]  ( .D(n5566), .CK(CLK), .QN(n7905) );
  DFF_X1 \REGISTERS_reg[23][49]  ( .D(n5565), .CK(CLK), .QN(n7908) );
  DFF_X1 \REGISTERS_reg[23][48]  ( .D(n5564), .CK(CLK), .QN(n7911) );
  DFF_X1 \REGISTERS_reg[23][47]  ( .D(n5563), .CK(CLK), .QN(n7914) );
  DFF_X1 \REGISTERS_reg[23][46]  ( .D(n5562), .CK(CLK), .QN(n7917) );
  DFF_X1 \REGISTERS_reg[23][45]  ( .D(n5561), .CK(CLK), .QN(n7920) );
  DFF_X1 \REGISTERS_reg[23][44]  ( .D(n5560), .CK(CLK), .QN(n7923) );
  DFF_X1 \REGISTERS_reg[23][43]  ( .D(n5559), .CK(CLK), .QN(n7926) );
  DFF_X1 \REGISTERS_reg[23][42]  ( .D(n5558), .CK(CLK), .QN(n7929) );
  DFF_X1 \REGISTERS_reg[23][41]  ( .D(n5557), .CK(CLK), .QN(n7932) );
  DFF_X1 \REGISTERS_reg[23][40]  ( .D(n5556), .CK(CLK), .QN(n7935) );
  DFF_X1 \REGISTERS_reg[23][39]  ( .D(n5555), .CK(CLK), .QN(n7938) );
  DFF_X1 \REGISTERS_reg[23][38]  ( .D(n5554), .CK(CLK), .QN(n7941) );
  DFF_X1 \REGISTERS_reg[23][37]  ( .D(n5553), .CK(CLK), .QN(n7944) );
  DFF_X1 \REGISTERS_reg[23][36]  ( .D(n5552), .CK(CLK), .QN(n7947) );
  DFF_X1 \REGISTERS_reg[23][35]  ( .D(n5551), .CK(CLK), .QN(n7950) );
  DFF_X1 \REGISTERS_reg[23][34]  ( .D(n5550), .CK(CLK), .QN(n7953) );
  DFF_X1 \REGISTERS_reg[23][33]  ( .D(n5549), .CK(CLK), .QN(n7956) );
  DFF_X1 \REGISTERS_reg[23][32]  ( .D(n5548), .CK(CLK), .QN(n7959) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n5547), .CK(CLK), .QN(n7962) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n5546), .CK(CLK), .QN(n7965) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n5545), .CK(CLK), .QN(n7968) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n5544), .CK(CLK), .QN(n7971) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n5543), .CK(CLK), .QN(n7974) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n5542), .CK(CLK), .QN(n7977) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n5541), .CK(CLK), .QN(n7980) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n5540), .CK(CLK), .QN(n7983) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n5539), .CK(CLK), .QN(n7986) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n5538), .CK(CLK), .QN(n7989) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n5537), .CK(CLK), .QN(n7992) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n5536), .CK(CLK), .QN(n7995) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n5535), .CK(CLK), .QN(n7998) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n5534), .CK(CLK), .QN(n8001) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n5533), .CK(CLK), .QN(n8004) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n5532), .CK(CLK), .QN(n8007) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n5531), .CK(CLK), .QN(n8010) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n5530), .CK(CLK), .QN(n8013) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n5529), .CK(CLK), .QN(n8016) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n5528), .CK(CLK), .QN(n8019) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n5527), .CK(CLK), .QN(n8022) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n5526), .CK(CLK), .QN(n8025) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n5525), .CK(CLK), .QN(n8028) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n5524), .CK(CLK), .QN(n8031) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n5523), .CK(CLK), .QN(n8034) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n5522), .CK(CLK), .QN(n8037) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n5521), .CK(CLK), .QN(n8040) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n5520), .CK(CLK), .QN(n8043) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n5519), .CK(CLK), .QN(n8046) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n5518), .CK(CLK), .QN(n8049) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n5517), .CK(CLK), .QN(n8052) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n5516), .CK(CLK), .QN(n8055) );
  DFF_X1 \REGISTERS_reg[29][62]  ( .D(n5194), .CK(CLK), .QN(n7739) );
  DFF_X1 \REGISTERS_reg[29][61]  ( .D(n5193), .CK(CLK), .QN(n7741) );
  DFF_X1 \REGISTERS_reg[29][60]  ( .D(n5192), .CK(CLK), .QN(n7743) );
  DFF_X1 \REGISTERS_reg[29][59]  ( .D(n5191), .CK(CLK), .QN(n7745) );
  DFF_X1 \REGISTERS_reg[29][58]  ( .D(n5190), .CK(CLK), .QN(n7747) );
  DFF_X1 \REGISTERS_reg[29][57]  ( .D(n5189), .CK(CLK), .QN(n7749) );
  DFF_X1 \REGISTERS_reg[29][56]  ( .D(n5188), .CK(CLK), .QN(n7751) );
  DFF_X1 \REGISTERS_reg[29][55]  ( .D(n5187), .CK(CLK), .QN(n7753) );
  DFF_X1 \REGISTERS_reg[29][54]  ( .D(n5186), .CK(CLK), .QN(n7755) );
  DFF_X1 \REGISTERS_reg[29][53]  ( .D(n5185), .CK(CLK), .QN(n7757) );
  DFF_X1 \REGISTERS_reg[29][52]  ( .D(n5184), .CK(CLK), .QN(n7759) );
  DFF_X1 \REGISTERS_reg[29][51]  ( .D(n5183), .CK(CLK), .QN(n7761) );
  DFF_X1 \REGISTERS_reg[29][50]  ( .D(n5182), .CK(CLK), .QN(n7763) );
  DFF_X1 \REGISTERS_reg[29][49]  ( .D(n5181), .CK(CLK), .QN(n7765) );
  DFF_X1 \REGISTERS_reg[29][48]  ( .D(n5180), .CK(CLK), .QN(n7767) );
  DFF_X1 \REGISTERS_reg[29][47]  ( .D(n5179), .CK(CLK), .QN(n7769) );
  DFF_X1 \REGISTERS_reg[29][46]  ( .D(n5178), .CK(CLK), .QN(n7771) );
  DFF_X1 \REGISTERS_reg[29][45]  ( .D(n5177), .CK(CLK), .QN(n7773) );
  DFF_X1 \REGISTERS_reg[29][44]  ( .D(n5176), .CK(CLK), .QN(n7775) );
  DFF_X1 \REGISTERS_reg[29][43]  ( .D(n5175), .CK(CLK), .QN(n7777) );
  DFF_X1 \REGISTERS_reg[29][42]  ( .D(n5174), .CK(CLK), .QN(n7779) );
  DFF_X1 \REGISTERS_reg[29][41]  ( .D(n5173), .CK(CLK), .QN(n7781) );
  DFF_X1 \REGISTERS_reg[29][40]  ( .D(n5172), .CK(CLK), .QN(n7783) );
  DFF_X1 \REGISTERS_reg[29][39]  ( .D(n5171), .CK(CLK), .QN(n7785) );
  DFF_X1 \REGISTERS_reg[29][38]  ( .D(n5170), .CK(CLK), .QN(n7787) );
  DFF_X1 \REGISTERS_reg[29][37]  ( .D(n5169), .CK(CLK), .QN(n7789) );
  DFF_X1 \REGISTERS_reg[29][36]  ( .D(n5168), .CK(CLK), .QN(n7791) );
  DFF_X1 \REGISTERS_reg[29][35]  ( .D(n5167), .CK(CLK), .QN(n7793) );
  DFF_X1 \REGISTERS_reg[29][34]  ( .D(n5166), .CK(CLK), .QN(n7795) );
  DFF_X1 \REGISTERS_reg[29][33]  ( .D(n5165), .CK(CLK), .QN(n7797) );
  DFF_X1 \REGISTERS_reg[29][32]  ( .D(n5164), .CK(CLK), .QN(n7799) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n5163), .CK(CLK), .QN(n7801) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n5162), .CK(CLK), .QN(n7803) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n5161), .CK(CLK), .QN(n7805) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n5160), .CK(CLK), .QN(n7807) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n5159), .CK(CLK), .QN(n7809) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n5158), .CK(CLK), .QN(n7811) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n5157), .CK(CLK), .QN(n7813) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n5156), .CK(CLK), .QN(n7815) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n5155), .CK(CLK), .QN(n7817) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n5154), .CK(CLK), .QN(n7819) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n5153), .CK(CLK), .QN(n7821) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n5152), .CK(CLK), .QN(n7823) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n5151), .CK(CLK), .QN(n7825) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n5150), .CK(CLK), .QN(n7827) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n5149), .CK(CLK), .QN(n7829) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n5148), .CK(CLK), .QN(n7831) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n5147), .CK(CLK), .QN(n7833) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n5146), .CK(CLK), .QN(n7835) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n5145), .CK(CLK), .QN(n7837) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n5144), .CK(CLK), .QN(n7839) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n5143), .CK(CLK), .QN(n7841) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n5142), .CK(CLK), .QN(n7843) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n5141), .CK(CLK), .QN(n7845) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n5140), .CK(CLK), .QN(n7847) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n5139), .CK(CLK), .QN(n7849) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n5138), .CK(CLK), .QN(n7851) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n5137), .CK(CLK), .QN(n7853) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n5136), .CK(CLK), .QN(n7855) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n5135), .CK(CLK), .QN(n7857) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n5134), .CK(CLK), .QN(n7859) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n5133), .CK(CLK), .QN(n7861) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n5132), .CK(CLK), .QN(n7863) );
  DFF_X1 \OUT1_reg[59]  ( .D(n4999), .CK(CLK), .Q(OUT1[59]) );
  DFF_X1 \OUT1_reg[58]  ( .D(n4998), .CK(CLK), .Q(OUT1[58]) );
  DFF_X1 \OUT1_reg[57]  ( .D(n4997), .CK(CLK), .Q(OUT1[57]) );
  DFF_X1 \OUT1_reg[56]  ( .D(n4996), .CK(CLK), .Q(OUT1[56]) );
  DFF_X1 \OUT1_reg[55]  ( .D(n4995), .CK(CLK), .Q(OUT1[55]) );
  DFF_X1 \OUT1_reg[54]  ( .D(n4994), .CK(CLK), .Q(OUT1[54]) );
  DFF_X1 \OUT1_reg[53]  ( .D(n4993), .CK(CLK), .Q(OUT1[53]) );
  DFF_X1 \OUT1_reg[52]  ( .D(n4992), .CK(CLK), .Q(OUT1[52]) );
  DFF_X1 \OUT1_reg[51]  ( .D(n4991), .CK(CLK), .Q(OUT1[51]) );
  DFF_X1 \OUT1_reg[50]  ( .D(n4990), .CK(CLK), .Q(OUT1[50]) );
  DFF_X1 \OUT1_reg[49]  ( .D(n4989), .CK(CLK), .Q(OUT1[49]) );
  DFF_X1 \OUT1_reg[48]  ( .D(n4988), .CK(CLK), .Q(OUT1[48]) );
  DFF_X1 \OUT1_reg[47]  ( .D(n4987), .CK(CLK), .Q(OUT1[47]) );
  DFF_X1 \OUT1_reg[46]  ( .D(n4986), .CK(CLK), .Q(OUT1[46]) );
  DFF_X1 \OUT1_reg[45]  ( .D(n4985), .CK(CLK), .Q(OUT1[45]) );
  DFF_X1 \OUT1_reg[44]  ( .D(n4984), .CK(CLK), .Q(OUT1[44]) );
  DFF_X1 \OUT1_reg[43]  ( .D(n4983), .CK(CLK), .Q(OUT1[43]) );
  DFF_X1 \OUT1_reg[42]  ( .D(n4982), .CK(CLK), .Q(OUT1[42]) );
  DFF_X1 \OUT1_reg[41]  ( .D(n4981), .CK(CLK), .Q(OUT1[41]) );
  DFF_X1 \OUT1_reg[40]  ( .D(n4980), .CK(CLK), .Q(OUT1[40]) );
  DFF_X1 \OUT1_reg[39]  ( .D(n4979), .CK(CLK), .Q(OUT1[39]) );
  DFF_X1 \OUT1_reg[38]  ( .D(n4978), .CK(CLK), .Q(OUT1[38]) );
  DFF_X1 \OUT1_reg[37]  ( .D(n4977), .CK(CLK), .Q(OUT1[37]) );
  DFF_X1 \OUT1_reg[36]  ( .D(n4976), .CK(CLK), .Q(OUT1[36]) );
  DFF_X1 \OUT1_reg[35]  ( .D(n4975), .CK(CLK), .Q(OUT1[35]) );
  DFF_X1 \OUT1_reg[34]  ( .D(n4974), .CK(CLK), .Q(OUT1[34]) );
  DFF_X1 \OUT1_reg[33]  ( .D(n4973), .CK(CLK), .Q(OUT1[33]) );
  DFF_X1 \OUT1_reg[32]  ( .D(n4972), .CK(CLK), .Q(OUT1[32]) );
  DFF_X1 \OUT1_reg[31]  ( .D(n4971), .CK(CLK), .Q(OUT1[31]) );
  DFF_X1 \OUT1_reg[30]  ( .D(n4970), .CK(CLK), .Q(OUT1[30]) );
  DFF_X1 \OUT1_reg[29]  ( .D(n4969), .CK(CLK), .Q(OUT1[29]) );
  DFF_X1 \OUT1_reg[28]  ( .D(n4968), .CK(CLK), .Q(OUT1[28]) );
  DFF_X1 \OUT1_reg[27]  ( .D(n4967), .CK(CLK), .Q(OUT1[27]) );
  DFF_X1 \OUT1_reg[26]  ( .D(n4966), .CK(CLK), .Q(OUT1[26]) );
  DFF_X1 \OUT1_reg[25]  ( .D(n4965), .CK(CLK), .Q(OUT1[25]) );
  DFF_X1 \OUT1_reg[24]  ( .D(n4964), .CK(CLK), .Q(OUT1[24]) );
  DFF_X1 \OUT1_reg[23]  ( .D(n4963), .CK(CLK), .Q(OUT1[23]) );
  DFF_X1 \OUT1_reg[22]  ( .D(n4962), .CK(CLK), .Q(OUT1[22]) );
  DFF_X1 \OUT1_reg[21]  ( .D(n4961), .CK(CLK), .Q(OUT1[21]) );
  DFF_X1 \OUT1_reg[20]  ( .D(n4960), .CK(CLK), .Q(OUT1[20]) );
  DFF_X1 \OUT1_reg[19]  ( .D(n4959), .CK(CLK), .Q(OUT1[19]) );
  DFF_X1 \OUT1_reg[18]  ( .D(n4958), .CK(CLK), .Q(OUT1[18]) );
  DFF_X1 \OUT1_reg[17]  ( .D(n4957), .CK(CLK), .Q(OUT1[17]) );
  DFF_X1 \OUT1_reg[16]  ( .D(n4956), .CK(CLK), .Q(OUT1[16]) );
  DFF_X1 \OUT1_reg[15]  ( .D(n4955), .CK(CLK), .Q(OUT1[15]) );
  DFF_X1 \OUT1_reg[14]  ( .D(n4954), .CK(CLK), .Q(OUT1[14]) );
  DFF_X1 \OUT1_reg[13]  ( .D(n4953), .CK(CLK), .Q(OUT1[13]) );
  DFF_X1 \OUT1_reg[12]  ( .D(n4952), .CK(CLK), .Q(OUT1[12]) );
  DFF_X1 \OUT1_reg[11]  ( .D(n4951), .CK(CLK), .Q(OUT1[11]) );
  DFF_X1 \OUT1_reg[10]  ( .D(n4950), .CK(CLK), .Q(OUT1[10]) );
  DFF_X1 \OUT1_reg[9]  ( .D(n4949), .CK(CLK), .Q(OUT1[9]) );
  DFF_X1 \OUT1_reg[8]  ( .D(n4948), .CK(CLK), .Q(OUT1[8]) );
  DFF_X1 \OUT1_reg[7]  ( .D(n4947), .CK(CLK), .Q(OUT1[7]) );
  DFF_X1 \OUT1_reg[6]  ( .D(n4946), .CK(CLK), .Q(OUT1[6]) );
  DFF_X1 \OUT1_reg[5]  ( .D(n4945), .CK(CLK), .Q(OUT1[5]) );
  DFF_X1 \OUT1_reg[4]  ( .D(n4944), .CK(CLK), .Q(OUT1[4]) );
  DFF_X1 \OUT1_reg[3]  ( .D(n4943), .CK(CLK), .Q(OUT1[3]) );
  DFF_X1 \OUT1_reg[2]  ( .D(n4942), .CK(CLK), .Q(OUT1[2]) );
  DFF_X1 \OUT1_reg[1]  ( .D(n4941), .CK(CLK), .Q(OUT1[1]) );
  DFF_X1 \OUT1_reg[0]  ( .D(n4940), .CK(CLK), .Q(OUT1[0]) );
  DFF_X1 \OUT2_reg[31]  ( .D(n4907), .CK(CLK), .Q(OUT2[31]) );
  DFF_X1 \OUT2_reg[30]  ( .D(n4906), .CK(CLK), .Q(OUT2[30]) );
  DFF_X1 \OUT2_reg[29]  ( .D(n4905), .CK(CLK), .Q(OUT2[29]) );
  DFF_X1 \OUT2_reg[28]  ( .D(n4904), .CK(CLK), .Q(OUT2[28]) );
  DFF_X1 \OUT2_reg[27]  ( .D(n4903), .CK(CLK), .Q(OUT2[27]) );
  DFF_X1 \OUT2_reg[26]  ( .D(n4902), .CK(CLK), .Q(OUT2[26]) );
  DFF_X1 \OUT2_reg[25]  ( .D(n4901), .CK(CLK), .Q(OUT2[25]) );
  DFF_X1 \OUT2_reg[24]  ( .D(n4900), .CK(CLK), .Q(OUT2[24]) );
  DFF_X1 \OUT2_reg[23]  ( .D(n4899), .CK(CLK), .Q(OUT2[23]) );
  DFF_X1 \OUT2_reg[22]  ( .D(n4898), .CK(CLK), .Q(OUT2[22]) );
  DFF_X1 \OUT2_reg[21]  ( .D(n4897), .CK(CLK), .Q(OUT2[21]) );
  DFF_X1 \OUT2_reg[20]  ( .D(n4896), .CK(CLK), .Q(OUT2[20]) );
  DFF_X1 \OUT2_reg[19]  ( .D(n4895), .CK(CLK), .Q(OUT2[19]) );
  DFF_X1 \OUT2_reg[18]  ( .D(n4894), .CK(CLK), .Q(OUT2[18]) );
  DFF_X1 \OUT2_reg[17]  ( .D(n4893), .CK(CLK), .Q(OUT2[17]) );
  DFF_X1 \OUT2_reg[16]  ( .D(n4892), .CK(CLK), .Q(OUT2[16]) );
  DFF_X1 \OUT2_reg[15]  ( .D(n4891), .CK(CLK), .Q(OUT2[15]) );
  DFF_X1 \OUT2_reg[14]  ( .D(n4890), .CK(CLK), .Q(OUT2[14]) );
  DFF_X1 \OUT2_reg[13]  ( .D(n4889), .CK(CLK), .Q(OUT2[13]) );
  DFF_X1 \OUT2_reg[12]  ( .D(n4888), .CK(CLK), .Q(OUT2[12]) );
  DFF_X1 \OUT2_reg[11]  ( .D(n4887), .CK(CLK), .Q(OUT2[11]) );
  DFF_X1 \OUT2_reg[10]  ( .D(n4886), .CK(CLK), .Q(OUT2[10]) );
  DFF_X1 \OUT2_reg[9]  ( .D(n4885), .CK(CLK), .Q(OUT2[9]) );
  DFF_X1 \OUT2_reg[8]  ( .D(n4884), .CK(CLK), .Q(OUT2[8]) );
  DFF_X1 \OUT2_reg[7]  ( .D(n4883), .CK(CLK), .Q(OUT2[7]) );
  DFF_X1 \OUT2_reg[6]  ( .D(n4882), .CK(CLK), .Q(OUT2[6]) );
  DFF_X1 \OUT2_reg[5]  ( .D(n4881), .CK(CLK), .Q(OUT2[5]) );
  DFF_X1 \OUT2_reg[4]  ( .D(n4880), .CK(CLK), .Q(OUT2[4]) );
  DFF_X1 \OUT2_reg[3]  ( .D(n4879), .CK(CLK), .Q(OUT2[3]) );
  DFF_X1 \OUT2_reg[2]  ( .D(n4878), .CK(CLK), .Q(OUT2[2]) );
  DFF_X1 \OUT2_reg[1]  ( .D(n4877), .CK(CLK), .Q(OUT2[1]) );
  DFF_X1 \OUT2_reg[0]  ( .D(n4876), .CK(CLK), .Q(OUT2[0]) );
  NAND3_X1 U11147 ( .A1(n12184), .A2(n12183), .A3(n13652), .ZN(n13636) );
  NAND3_X1 U11148 ( .A1(n13652), .A2(n12183), .A3(ADD_WR[3]), .ZN(n13654) );
  NAND3_X1 U11149 ( .A1(n13652), .A2(n12184), .A3(ADD_WR[4]), .ZN(n13663) );
  NAND3_X1 U11150 ( .A1(n12186), .A2(n12185), .A3(n12187), .ZN(n13637) );
  NAND3_X1 U11151 ( .A1(n12186), .A2(n12185), .A3(ADD_WR[0]), .ZN(n13639) );
  NAND3_X1 U11152 ( .A1(n12187), .A2(n12185), .A3(ADD_WR[1]), .ZN(n13641) );
  NAND3_X1 U11153 ( .A1(ADD_WR[0]), .A2(n12185), .A3(ADD_WR[1]), .ZN(n13643)
         );
  NAND3_X1 U11154 ( .A1(n12187), .A2(n12186), .A3(ADD_WR[2]), .ZN(n13645) );
  NAND3_X1 U11155 ( .A1(ADD_WR[0]), .A2(n12186), .A3(ADD_WR[2]), .ZN(n13647)
         );
  NAND3_X1 U11156 ( .A1(ADD_WR[1]), .A2(n12187), .A3(ADD_WR[2]), .ZN(n13649)
         );
  NAND3_X1 U11157 ( .A1(ADD_WR[3]), .A2(n13652), .A3(ADD_WR[4]), .ZN(n13672)
         );
  NAND3_X1 U11158 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n13651) );
  NAND3_X1 U11159 ( .A1(n14857), .A2(n16685), .A3(n14860), .ZN(n13687) );
  NAND3_X1 U11160 ( .A1(n14856), .A2(n14861), .A3(n14862), .ZN(n13686) );
  NAND3_X1 U11161 ( .A1(n14865), .A2(n16686), .A3(n14860), .ZN(n13692) );
  NAND3_X1 U11162 ( .A1(n14865), .A2(n16686), .A3(n14866), .ZN(n13691) );
  NAND3_X1 U11163 ( .A1(n14862), .A2(n16686), .A3(n14859), .ZN(n13697) );
  NAND3_X1 U11164 ( .A1(n14857), .A2(n16686), .A3(n14859), .ZN(n13696) );
  NAND3_X1 U11165 ( .A1(n16686), .A2(n14861), .A3(n14865), .ZN(n13702) );
  NAND3_X1 U11166 ( .A1(n14864), .A2(n16686), .A3(n14857), .ZN(n13701) );
  NAND3_X1 U11167 ( .A1(n14862), .A2(n16685), .A3(n14866), .ZN(n13722) );
  NAND3_X1 U11168 ( .A1(n14862), .A2(n16685), .A3(n14855), .ZN(n13721) );
  NAND3_X1 U11169 ( .A1(n14862), .A2(n16685), .A3(n14860), .ZN(n13727) );
  NAND3_X1 U11170 ( .A1(n14865), .A2(n16685), .A3(n14859), .ZN(n13726) );
  XOR2_X1 U11171 ( .A(ADD_WR[4]), .B(ADD_RD1[4]), .Z(n14886) );
  XOR2_X1 U11172 ( .A(ADD_WR[2]), .B(ADD_RD1[2]), .Z(n14885) );
  XOR2_X1 U11173 ( .A(n12192), .B(ADD_WR[0]), .Z(n14883) );
  XOR2_X1 U11174 ( .A(n12191), .B(ADD_WR[1]), .Z(n14882) );
  XOR2_X1 U11175 ( .A(n12184), .B(ADD_RD1[3]), .Z(n14881) );
  NAND3_X1 U11176 ( .A1(n16065), .A2(n16480), .A3(n16068), .ZN(n14895) );
  NAND3_X1 U11177 ( .A1(n16064), .A2(n16069), .A3(n16070), .ZN(n14894) );
  NAND3_X1 U11178 ( .A1(n16073), .A2(n16481), .A3(n16068), .ZN(n14900) );
  NAND3_X1 U11179 ( .A1(n16073), .A2(n16481), .A3(n16074), .ZN(n14899) );
  NAND3_X1 U11180 ( .A1(n16070), .A2(n16481), .A3(n16067), .ZN(n14905) );
  NAND3_X1 U11181 ( .A1(n16065), .A2(n16481), .A3(n16067), .ZN(n14904) );
  NAND3_X1 U11182 ( .A1(n16481), .A2(n16069), .A3(n16073), .ZN(n14910) );
  NAND3_X1 U11183 ( .A1(n16072), .A2(n16481), .A3(n16065), .ZN(n14909) );
  NAND3_X1 U11184 ( .A1(n16070), .A2(n16480), .A3(n16074), .ZN(n14930) );
  NAND3_X1 U11185 ( .A1(n16070), .A2(n16480), .A3(n16063), .ZN(n14929) );
  NAND3_X1 U11186 ( .A1(n16070), .A2(n16480), .A3(n16068), .ZN(n14935) );
  NAND3_X1 U11187 ( .A1(n16073), .A2(n16480), .A3(n16067), .ZN(n14934) );
  XOR2_X1 U11188 ( .A(ADD_WR[4]), .B(ADD_RD2[4]), .Z(n16094) );
  XOR2_X1 U11189 ( .A(ADD_WR[2]), .B(ADD_RD2[2]), .Z(n16093) );
  XOR2_X1 U11190 ( .A(n12197), .B(ADD_WR[0]), .Z(n16091) );
  XOR2_X1 U11191 ( .A(n12196), .B(ADD_WR[1]), .Z(n16090) );
  XOR2_X1 U11192 ( .A(n12184), .B(ADD_RD2[3]), .Z(n16089) );
  DFF_X1 \REGISTERS_reg[28][63]  ( .D(n5259), .CK(CLK), .Q(n13379), .QN(n7609)
         );
  DFF_X1 \REGISTERS_reg[28][62]  ( .D(n5258), .CK(CLK), .Q(n13380), .QN(n7611)
         );
  DFF_X1 \REGISTERS_reg[28][61]  ( .D(n5257), .CK(CLK), .Q(n13381), .QN(n7613)
         );
  DFF_X1 \REGISTERS_reg[28][60]  ( .D(n5256), .CK(CLK), .Q(n13382), .QN(n7615)
         );
  DFF_X1 \REGISTERS_reg[25][63]  ( .D(n5451), .CK(CLK), .Q(n13187), .QN(n7244)
         );
  DFF_X1 \REGISTERS_reg[25][62]  ( .D(n5450), .CK(CLK), .Q(n13188), .QN(n7245)
         );
  DFF_X1 \REGISTERS_reg[25][61]  ( .D(n5449), .CK(CLK), .Q(n13189), .QN(n7246)
         );
  DFF_X1 \REGISTERS_reg[25][60]  ( .D(n5448), .CK(CLK), .Q(n13190), .QN(n7247)
         );
  DFF_X1 \REGISTERS_reg[24][63]  ( .D(n5515), .CK(CLK), .Q(n13123), .QN(n7867)
         );
  DFF_X1 \REGISTERS_reg[24][62]  ( .D(n5514), .CK(CLK), .Q(n13124), .QN(n7870)
         );
  DFF_X1 \REGISTERS_reg[24][61]  ( .D(n5513), .CK(CLK), .Q(n13125), .QN(n7873)
         );
  DFF_X1 \REGISTERS_reg[24][60]  ( .D(n5512), .CK(CLK), .Q(n13126), .QN(n7876)
         );
  DFF_X1 \REGISTERS_reg[22][63]  ( .D(n5643), .CK(CLK), .Q(n13059), .QN(n7309)
         );
  DFF_X1 \REGISTERS_reg[22][62]  ( .D(n5642), .CK(CLK), .Q(n13060), .QN(n7311)
         );
  DFF_X1 \REGISTERS_reg[22][61]  ( .D(n5641), .CK(CLK), .Q(n13061), .QN(n7313)
         );
  DFF_X1 \REGISTERS_reg[22][60]  ( .D(n5640), .CK(CLK), .Q(n13062), .QN(n7315)
         );
  DFF_X1 \REGISTERS_reg[5][63]  ( .D(n6731), .CK(CLK), .Q(n12390), .QN(n7052)
         );
  DFF_X1 \REGISTERS_reg[5][62]  ( .D(n6730), .CK(CLK), .Q(n12391), .QN(n7053)
         );
  DFF_X1 \REGISTERS_reg[5][61]  ( .D(n6729), .CK(CLK), .Q(n12392), .QN(n7054)
         );
  DFF_X1 \REGISTERS_reg[5][60]  ( .D(n6728), .CK(CLK), .Q(n12393), .QN(n7055)
         );
  DFF_X1 \REGISTERS_reg[4][63]  ( .D(n6795), .CK(CLK), .Q(n12326), .QN(n16100)
         );
  DFF_X1 \REGISTERS_reg[4][62]  ( .D(n6794), .CK(CLK), .Q(n12327), .QN(n16105)
         );
  DFF_X1 \REGISTERS_reg[4][61]  ( .D(n6793), .CK(CLK), .Q(n12328), .QN(n16110)
         );
  DFF_X1 \REGISTERS_reg[4][60]  ( .D(n6792), .CK(CLK), .Q(n12329), .QN(n16115)
         );
  DFF_X1 \REGISTERS_reg[1][63]  ( .D(n6987), .CK(CLK), .Q(n12262), .QN(n7865)
         );
  DFF_X1 \REGISTERS_reg[1][62]  ( .D(n6986), .CK(CLK), .Q(n12263), .QN(n7868)
         );
  DFF_X1 \REGISTERS_reg[1][61]  ( .D(n6985), .CK(CLK), .Q(n12264), .QN(n7871)
         );
  DFF_X1 \REGISTERS_reg[1][60]  ( .D(n6984), .CK(CLK), .Q(n12265), .QN(n7874)
         );
  DFF_X1 \REGISTERS_reg[0][63]  ( .D(n7051), .CK(CLK), .Q(n12198), .QN(n7308)
         );
  DFF_X1 \REGISTERS_reg[0][62]  ( .D(n7050), .CK(CLK), .Q(n12199), .QN(n7310)
         );
  DFF_X1 \REGISTERS_reg[0][61]  ( .D(n7049), .CK(CLK), .Q(n12200), .QN(n7312)
         );
  DFF_X1 \REGISTERS_reg[0][60]  ( .D(n7048), .CK(CLK), .Q(n12201), .QN(n7314)
         );
  DFF_X1 \REGISTERS_reg[28][59]  ( .D(n5255), .CK(CLK), .Q(n13383), .QN(n7617)
         );
  DFF_X1 \REGISTERS_reg[28][58]  ( .D(n5254), .CK(CLK), .Q(n13384), .QN(n7619)
         );
  DFF_X1 \REGISTERS_reg[28][57]  ( .D(n5253), .CK(CLK), .Q(n13385), .QN(n7621)
         );
  DFF_X1 \REGISTERS_reg[28][56]  ( .D(n5252), .CK(CLK), .Q(n13386), .QN(n7623)
         );
  DFF_X1 \REGISTERS_reg[28][55]  ( .D(n5251), .CK(CLK), .Q(n13387), .QN(n7625)
         );
  DFF_X1 \REGISTERS_reg[28][54]  ( .D(n5250), .CK(CLK), .Q(n13388), .QN(n7627)
         );
  DFF_X1 \REGISTERS_reg[28][53]  ( .D(n5249), .CK(CLK), .Q(n13389), .QN(n7629)
         );
  DFF_X1 \REGISTERS_reg[28][52]  ( .D(n5248), .CK(CLK), .Q(n13390), .QN(n7631)
         );
  DFF_X1 \REGISTERS_reg[28][51]  ( .D(n5247), .CK(CLK), .Q(n13391), .QN(n7633)
         );
  DFF_X1 \REGISTERS_reg[28][50]  ( .D(n5246), .CK(CLK), .Q(n13392), .QN(n7635)
         );
  DFF_X1 \REGISTERS_reg[28][49]  ( .D(n5245), .CK(CLK), .Q(n13393), .QN(n7637)
         );
  DFF_X1 \REGISTERS_reg[28][48]  ( .D(n5244), .CK(CLK), .Q(n13394), .QN(n7639)
         );
  DFF_X1 \REGISTERS_reg[28][47]  ( .D(n5243), .CK(CLK), .Q(n13395), .QN(n7641)
         );
  DFF_X1 \REGISTERS_reg[28][46]  ( .D(n5242), .CK(CLK), .Q(n13396), .QN(n7643)
         );
  DFF_X1 \REGISTERS_reg[28][45]  ( .D(n5241), .CK(CLK), .Q(n13397), .QN(n7645)
         );
  DFF_X1 \REGISTERS_reg[28][44]  ( .D(n5240), .CK(CLK), .Q(n13398), .QN(n7647)
         );
  DFF_X1 \REGISTERS_reg[28][43]  ( .D(n5239), .CK(CLK), .Q(n13399), .QN(n7649)
         );
  DFF_X1 \REGISTERS_reg[28][42]  ( .D(n5238), .CK(CLK), .Q(n13400), .QN(n7651)
         );
  DFF_X1 \REGISTERS_reg[28][41]  ( .D(n5237), .CK(CLK), .Q(n13401), .QN(n7653)
         );
  DFF_X1 \REGISTERS_reg[28][40]  ( .D(n5236), .CK(CLK), .Q(n13402), .QN(n7655)
         );
  DFF_X1 \REGISTERS_reg[28][39]  ( .D(n5235), .CK(CLK), .Q(n13403), .QN(n7657)
         );
  DFF_X1 \REGISTERS_reg[28][38]  ( .D(n5234), .CK(CLK), .Q(n13404), .QN(n7659)
         );
  DFF_X1 \REGISTERS_reg[28][37]  ( .D(n5233), .CK(CLK), .Q(n13405), .QN(n7661)
         );
  DFF_X1 \REGISTERS_reg[28][36]  ( .D(n5232), .CK(CLK), .Q(n13406), .QN(n7663)
         );
  DFF_X1 \REGISTERS_reg[28][35]  ( .D(n5231), .CK(CLK), .Q(n13407), .QN(n7665)
         );
  DFF_X1 \REGISTERS_reg[28][34]  ( .D(n5230), .CK(CLK), .Q(n13408), .QN(n7667)
         );
  DFF_X1 \REGISTERS_reg[28][33]  ( .D(n5229), .CK(CLK), .Q(n13409), .QN(n7669)
         );
  DFF_X1 \REGISTERS_reg[28][32]  ( .D(n5228), .CK(CLK), .Q(n13410), .QN(n7671)
         );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n5227), .CK(CLK), .Q(n13411), .QN(n7673)
         );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n5226), .CK(CLK), .Q(n13412), .QN(n7675)
         );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n5225), .CK(CLK), .Q(n13413), .QN(n7677)
         );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n5224), .CK(CLK), .Q(n13414), .QN(n7679)
         );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n5223), .CK(CLK), .Q(n13415), .QN(n7681)
         );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n5222), .CK(CLK), .Q(n13416), .QN(n7683)
         );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n5221), .CK(CLK), .Q(n13417), .QN(n7685)
         );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n5220), .CK(CLK), .Q(n13418), .QN(n7687)
         );
  DFF_X1 \REGISTERS_reg[25][59]  ( .D(n5447), .CK(CLK), .Q(n13191), .QN(n7248)
         );
  DFF_X1 \REGISTERS_reg[25][58]  ( .D(n5446), .CK(CLK), .Q(n13192), .QN(n7249)
         );
  DFF_X1 \REGISTERS_reg[25][57]  ( .D(n5445), .CK(CLK), .Q(n13193), .QN(n7250)
         );
  DFF_X1 \REGISTERS_reg[25][56]  ( .D(n5444), .CK(CLK), .Q(n13194), .QN(n7251)
         );
  DFF_X1 \REGISTERS_reg[25][55]  ( .D(n5443), .CK(CLK), .Q(n13195), .QN(n7252)
         );
  DFF_X1 \REGISTERS_reg[25][54]  ( .D(n5442), .CK(CLK), .Q(n13196), .QN(n7253)
         );
  DFF_X1 \REGISTERS_reg[25][53]  ( .D(n5441), .CK(CLK), .Q(n13197), .QN(n7254)
         );
  DFF_X1 \REGISTERS_reg[25][52]  ( .D(n5440), .CK(CLK), .Q(n13198), .QN(n7255)
         );
  DFF_X1 \REGISTERS_reg[25][51]  ( .D(n5439), .CK(CLK), .Q(n13199), .QN(n7256)
         );
  DFF_X1 \REGISTERS_reg[25][50]  ( .D(n5438), .CK(CLK), .Q(n13200), .QN(n7257)
         );
  DFF_X1 \REGISTERS_reg[25][49]  ( .D(n5437), .CK(CLK), .Q(n13201), .QN(n7258)
         );
  DFF_X1 \REGISTERS_reg[25][48]  ( .D(n5436), .CK(CLK), .Q(n13202), .QN(n7259)
         );
  DFF_X1 \REGISTERS_reg[25][47]  ( .D(n5435), .CK(CLK), .Q(n13203), .QN(n7260)
         );
  DFF_X1 \REGISTERS_reg[25][46]  ( .D(n5434), .CK(CLK), .Q(n13204), .QN(n7261)
         );
  DFF_X1 \REGISTERS_reg[25][45]  ( .D(n5433), .CK(CLK), .Q(n13205), .QN(n7262)
         );
  DFF_X1 \REGISTERS_reg[25][44]  ( .D(n5432), .CK(CLK), .Q(n13206), .QN(n7263)
         );
  DFF_X1 \REGISTERS_reg[25][43]  ( .D(n5431), .CK(CLK), .Q(n13207), .QN(n7264)
         );
  DFF_X1 \REGISTERS_reg[25][42]  ( .D(n5430), .CK(CLK), .Q(n13208), .QN(n7265)
         );
  DFF_X1 \REGISTERS_reg[25][41]  ( .D(n5429), .CK(CLK), .Q(n13209), .QN(n7266)
         );
  DFF_X1 \REGISTERS_reg[25][40]  ( .D(n5428), .CK(CLK), .Q(n13210), .QN(n7267)
         );
  DFF_X1 \REGISTERS_reg[25][39]  ( .D(n5427), .CK(CLK), .Q(n13211), .QN(n7268)
         );
  DFF_X1 \REGISTERS_reg[25][38]  ( .D(n5426), .CK(CLK), .Q(n13212), .QN(n7269)
         );
  DFF_X1 \REGISTERS_reg[25][37]  ( .D(n5425), .CK(CLK), .Q(n13213), .QN(n7270)
         );
  DFF_X1 \REGISTERS_reg[25][36]  ( .D(n5424), .CK(CLK), .Q(n13214), .QN(n7271)
         );
  DFF_X1 \REGISTERS_reg[25][35]  ( .D(n5423), .CK(CLK), .Q(n13215), .QN(n7272)
         );
  DFF_X1 \REGISTERS_reg[25][34]  ( .D(n5422), .CK(CLK), .Q(n13216), .QN(n7273)
         );
  DFF_X1 \REGISTERS_reg[25][33]  ( .D(n5421), .CK(CLK), .Q(n13217), .QN(n7274)
         );
  DFF_X1 \REGISTERS_reg[25][32]  ( .D(n5420), .CK(CLK), .Q(n13218), .QN(n7275)
         );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n5419), .CK(CLK), .Q(n13219), .QN(n7276)
         );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n5418), .CK(CLK), .Q(n13220), .QN(n7277)
         );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n5417), .CK(CLK), .Q(n13221), .QN(n7278)
         );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n5416), .CK(CLK), .Q(n13222), .QN(n7279)
         );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n5415), .CK(CLK), .Q(n13223), .QN(n7280)
         );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n5414), .CK(CLK), .Q(n13224), .QN(n7281)
         );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n5413), .CK(CLK), .Q(n13225), .QN(n7282)
         );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n5412), .CK(CLK), .Q(n13226), .QN(n7283)
         );
  DFF_X1 \REGISTERS_reg[24][59]  ( .D(n5511), .CK(CLK), .Q(n13127), .QN(n7879)
         );
  DFF_X1 \REGISTERS_reg[24][58]  ( .D(n5510), .CK(CLK), .Q(n13128), .QN(n7882)
         );
  DFF_X1 \REGISTERS_reg[24][57]  ( .D(n5509), .CK(CLK), .Q(n13129), .QN(n7885)
         );
  DFF_X1 \REGISTERS_reg[24][56]  ( .D(n5508), .CK(CLK), .Q(n13130), .QN(n7888)
         );
  DFF_X1 \REGISTERS_reg[24][55]  ( .D(n5507), .CK(CLK), .Q(n13131), .QN(n7891)
         );
  DFF_X1 \REGISTERS_reg[24][54]  ( .D(n5506), .CK(CLK), .Q(n13132), .QN(n7894)
         );
  DFF_X1 \REGISTERS_reg[24][53]  ( .D(n5505), .CK(CLK), .Q(n13133), .QN(n7897)
         );
  DFF_X1 \REGISTERS_reg[24][52]  ( .D(n5504), .CK(CLK), .Q(n13134), .QN(n7900)
         );
  DFF_X1 \REGISTERS_reg[24][51]  ( .D(n5503), .CK(CLK), .Q(n13135), .QN(n7903)
         );
  DFF_X1 \REGISTERS_reg[24][50]  ( .D(n5502), .CK(CLK), .Q(n13136), .QN(n7906)
         );
  DFF_X1 \REGISTERS_reg[24][49]  ( .D(n5501), .CK(CLK), .Q(n13137), .QN(n7909)
         );
  DFF_X1 \REGISTERS_reg[24][48]  ( .D(n5500), .CK(CLK), .Q(n13138), .QN(n7912)
         );
  DFF_X1 \REGISTERS_reg[24][47]  ( .D(n5499), .CK(CLK), .Q(n13139), .QN(n7915)
         );
  DFF_X1 \REGISTERS_reg[24][46]  ( .D(n5498), .CK(CLK), .Q(n13140), .QN(n7918)
         );
  DFF_X1 \REGISTERS_reg[24][45]  ( .D(n5497), .CK(CLK), .Q(n13141), .QN(n7921)
         );
  DFF_X1 \REGISTERS_reg[24][44]  ( .D(n5496), .CK(CLK), .Q(n13142), .QN(n7924)
         );
  DFF_X1 \REGISTERS_reg[24][43]  ( .D(n5495), .CK(CLK), .Q(n13143), .QN(n7927)
         );
  DFF_X1 \REGISTERS_reg[24][42]  ( .D(n5494), .CK(CLK), .Q(n13144), .QN(n7930)
         );
  DFF_X1 \REGISTERS_reg[24][41]  ( .D(n5493), .CK(CLK), .Q(n13145), .QN(n7933)
         );
  DFF_X1 \REGISTERS_reg[24][40]  ( .D(n5492), .CK(CLK), .Q(n13146), .QN(n7936)
         );
  DFF_X1 \REGISTERS_reg[24][39]  ( .D(n5491), .CK(CLK), .Q(n13147), .QN(n7939)
         );
  DFF_X1 \REGISTERS_reg[24][38]  ( .D(n5490), .CK(CLK), .Q(n13148), .QN(n7942)
         );
  DFF_X1 \REGISTERS_reg[24][37]  ( .D(n5489), .CK(CLK), .Q(n13149), .QN(n7945)
         );
  DFF_X1 \REGISTERS_reg[24][36]  ( .D(n5488), .CK(CLK), .Q(n13150), .QN(n7948)
         );
  DFF_X1 \REGISTERS_reg[24][35]  ( .D(n5487), .CK(CLK), .Q(n13151), .QN(n7951)
         );
  DFF_X1 \REGISTERS_reg[24][34]  ( .D(n5486), .CK(CLK), .Q(n13152), .QN(n7954)
         );
  DFF_X1 \REGISTERS_reg[24][33]  ( .D(n5485), .CK(CLK), .Q(n13153), .QN(n7957)
         );
  DFF_X1 \REGISTERS_reg[24][32]  ( .D(n5484), .CK(CLK), .Q(n13154), .QN(n7960)
         );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n5483), .CK(CLK), .Q(n13155), .QN(n7963)
         );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n5482), .CK(CLK), .Q(n13156), .QN(n7966)
         );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n5481), .CK(CLK), .Q(n13157), .QN(n7969)
         );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n5480), .CK(CLK), .Q(n13158), .QN(n7972)
         );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n5479), .CK(CLK), .Q(n13159), .QN(n7975)
         );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n5478), .CK(CLK), .Q(n13160), .QN(n7978)
         );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n5477), .CK(CLK), .Q(n13161), .QN(n7981)
         );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n5476), .CK(CLK), .Q(n13162), .QN(n7984)
         );
  DFF_X1 \REGISTERS_reg[22][59]  ( .D(n5639), .CK(CLK), .Q(n13063), .QN(n7317)
         );
  DFF_X1 \REGISTERS_reg[22][58]  ( .D(n5638), .CK(CLK), .Q(n13064), .QN(n7319)
         );
  DFF_X1 \REGISTERS_reg[22][57]  ( .D(n5637), .CK(CLK), .Q(n13065), .QN(n7321)
         );
  DFF_X1 \REGISTERS_reg[22][56]  ( .D(n5636), .CK(CLK), .Q(n13066), .QN(n7323)
         );
  DFF_X1 \REGISTERS_reg[22][55]  ( .D(n5635), .CK(CLK), .Q(n13067), .QN(n7325)
         );
  DFF_X1 \REGISTERS_reg[22][54]  ( .D(n5634), .CK(CLK), .Q(n13068), .QN(n7327)
         );
  DFF_X1 \REGISTERS_reg[22][53]  ( .D(n5633), .CK(CLK), .Q(n13069), .QN(n7329)
         );
  DFF_X1 \REGISTERS_reg[22][52]  ( .D(n5632), .CK(CLK), .Q(n13070), .QN(n7331)
         );
  DFF_X1 \REGISTERS_reg[22][51]  ( .D(n5631), .CK(CLK), .Q(n13071), .QN(n7333)
         );
  DFF_X1 \REGISTERS_reg[22][50]  ( .D(n5630), .CK(CLK), .Q(n13072), .QN(n7335)
         );
  DFF_X1 \REGISTERS_reg[22][49]  ( .D(n5629), .CK(CLK), .Q(n13073), .QN(n7337)
         );
  DFF_X1 \REGISTERS_reg[22][48]  ( .D(n5628), .CK(CLK), .Q(n13074), .QN(n7339)
         );
  DFF_X1 \REGISTERS_reg[22][47]  ( .D(n5627), .CK(CLK), .Q(n13075), .QN(n7341)
         );
  DFF_X1 \REGISTERS_reg[22][46]  ( .D(n5626), .CK(CLK), .Q(n13076), .QN(n7343)
         );
  DFF_X1 \REGISTERS_reg[22][45]  ( .D(n5625), .CK(CLK), .Q(n13077), .QN(n7345)
         );
  DFF_X1 \REGISTERS_reg[22][44]  ( .D(n5624), .CK(CLK), .Q(n13078), .QN(n7347)
         );
  DFF_X1 \REGISTERS_reg[22][43]  ( .D(n5623), .CK(CLK), .Q(n13079), .QN(n7349)
         );
  DFF_X1 \REGISTERS_reg[22][42]  ( .D(n5622), .CK(CLK), .Q(n13080), .QN(n7351)
         );
  DFF_X1 \REGISTERS_reg[22][41]  ( .D(n5621), .CK(CLK), .Q(n13081), .QN(n7353)
         );
  DFF_X1 \REGISTERS_reg[22][40]  ( .D(n5620), .CK(CLK), .Q(n13082), .QN(n7355)
         );
  DFF_X1 \REGISTERS_reg[22][39]  ( .D(n5619), .CK(CLK), .Q(n13083), .QN(n7357)
         );
  DFF_X1 \REGISTERS_reg[22][38]  ( .D(n5618), .CK(CLK), .Q(n13084), .QN(n7359)
         );
  DFF_X1 \REGISTERS_reg[22][37]  ( .D(n5617), .CK(CLK), .Q(n13085), .QN(n7361)
         );
  DFF_X1 \REGISTERS_reg[22][36]  ( .D(n5616), .CK(CLK), .Q(n13086), .QN(n7363)
         );
  DFF_X1 \REGISTERS_reg[22][35]  ( .D(n5615), .CK(CLK), .Q(n13087), .QN(n7365)
         );
  DFF_X1 \REGISTERS_reg[22][34]  ( .D(n5614), .CK(CLK), .Q(n13088), .QN(n7367)
         );
  DFF_X1 \REGISTERS_reg[22][33]  ( .D(n5613), .CK(CLK), .Q(n13089), .QN(n7369)
         );
  DFF_X1 \REGISTERS_reg[22][32]  ( .D(n5612), .CK(CLK), .Q(n13090), .QN(n7371)
         );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n5611), .CK(CLK), .Q(n13091), .QN(n7373)
         );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n5610), .CK(CLK), .Q(n13092), .QN(n7375)
         );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n5609), .CK(CLK), .Q(n13093), .QN(n7377)
         );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n5608), .CK(CLK), .Q(n13094), .QN(n7379)
         );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n5607), .CK(CLK), .Q(n13095), .QN(n7381)
         );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n5606), .CK(CLK), .Q(n13096), .QN(n7383)
         );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n5605), .CK(CLK), .Q(n13097), .QN(n7385)
         );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n5604), .CK(CLK), .Q(n13098), .QN(n7387)
         );
  DFF_X1 \REGISTERS_reg[5][59]  ( .D(n6727), .CK(CLK), .Q(n12394), .QN(n7056)
         );
  DFF_X1 \REGISTERS_reg[5][58]  ( .D(n6726), .CK(CLK), .Q(n12395), .QN(n7057)
         );
  DFF_X1 \REGISTERS_reg[5][57]  ( .D(n6725), .CK(CLK), .Q(n12396), .QN(n7058)
         );
  DFF_X1 \REGISTERS_reg[5][56]  ( .D(n6724), .CK(CLK), .Q(n12397), .QN(n7059)
         );
  DFF_X1 \REGISTERS_reg[5][55]  ( .D(n6723), .CK(CLK), .Q(n12398), .QN(n7060)
         );
  DFF_X1 \REGISTERS_reg[5][54]  ( .D(n6722), .CK(CLK), .Q(n12399), .QN(n7061)
         );
  DFF_X1 \REGISTERS_reg[5][53]  ( .D(n6721), .CK(CLK), .Q(n12400), .QN(n7062)
         );
  DFF_X1 \REGISTERS_reg[5][52]  ( .D(n6720), .CK(CLK), .Q(n12401), .QN(n7063)
         );
  DFF_X1 \REGISTERS_reg[5][51]  ( .D(n6719), .CK(CLK), .Q(n12402), .QN(n7064)
         );
  DFF_X1 \REGISTERS_reg[5][50]  ( .D(n6718), .CK(CLK), .Q(n12403), .QN(n7065)
         );
  DFF_X1 \REGISTERS_reg[5][49]  ( .D(n6717), .CK(CLK), .Q(n12404), .QN(n7066)
         );
  DFF_X1 \REGISTERS_reg[5][48]  ( .D(n6716), .CK(CLK), .Q(n12405), .QN(n7067)
         );
  DFF_X1 \REGISTERS_reg[5][47]  ( .D(n6715), .CK(CLK), .Q(n12406), .QN(n7068)
         );
  DFF_X1 \REGISTERS_reg[5][46]  ( .D(n6714), .CK(CLK), .Q(n12407), .QN(n7069)
         );
  DFF_X1 \REGISTERS_reg[5][45]  ( .D(n6713), .CK(CLK), .Q(n12408), .QN(n7070)
         );
  DFF_X1 \REGISTERS_reg[5][44]  ( .D(n6712), .CK(CLK), .Q(n12409), .QN(n7071)
         );
  DFF_X1 \REGISTERS_reg[5][43]  ( .D(n6711), .CK(CLK), .Q(n12410), .QN(n7072)
         );
  DFF_X1 \REGISTERS_reg[5][42]  ( .D(n6710), .CK(CLK), .Q(n12411), .QN(n7073)
         );
  DFF_X1 \REGISTERS_reg[5][41]  ( .D(n6709), .CK(CLK), .Q(n12412), .QN(n7074)
         );
  DFF_X1 \REGISTERS_reg[5][40]  ( .D(n6708), .CK(CLK), .Q(n12413), .QN(n7075)
         );
  DFF_X1 \REGISTERS_reg[5][39]  ( .D(n6707), .CK(CLK), .Q(n12414), .QN(n7076)
         );
  DFF_X1 \REGISTERS_reg[5][38]  ( .D(n6706), .CK(CLK), .Q(n12415), .QN(n7077)
         );
  DFF_X1 \REGISTERS_reg[5][37]  ( .D(n6705), .CK(CLK), .Q(n12416), .QN(n7078)
         );
  DFF_X1 \REGISTERS_reg[5][36]  ( .D(n6704), .CK(CLK), .Q(n12417), .QN(n7079)
         );
  DFF_X1 \REGISTERS_reg[5][35]  ( .D(n6703), .CK(CLK), .Q(n12418), .QN(n7080)
         );
  DFF_X1 \REGISTERS_reg[5][34]  ( .D(n6702), .CK(CLK), .Q(n12419), .QN(n7081)
         );
  DFF_X1 \REGISTERS_reg[5][33]  ( .D(n6701), .CK(CLK), .Q(n12420), .QN(n7082)
         );
  DFF_X1 \REGISTERS_reg[5][32]  ( .D(n6700), .CK(CLK), .Q(n12421), .QN(n7083)
         );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n6699), .CK(CLK), .Q(n12422), .QN(n7084)
         );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n6698), .CK(CLK), .Q(n12423), .QN(n7085)
         );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n6697), .CK(CLK), .Q(n12424), .QN(n7086)
         );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n6696), .CK(CLK), .Q(n12425), .QN(n7087)
         );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n6695), .CK(CLK), .Q(n12426), .QN(n7088)
         );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n6694), .CK(CLK), .Q(n12427), .QN(n7089)
         );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n6693), .CK(CLK), .Q(n12428), .QN(n7090)
         );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n6692), .CK(CLK), .Q(n12429), .QN(n7091)
         );
  DFF_X1 \REGISTERS_reg[4][59]  ( .D(n6791), .CK(CLK), .Q(n12330), .QN(n16120)
         );
  DFF_X1 \REGISTERS_reg[4][58]  ( .D(n6790), .CK(CLK), .Q(n12331), .QN(n16125)
         );
  DFF_X1 \REGISTERS_reg[4][57]  ( .D(n6789), .CK(CLK), .Q(n12332), .QN(n16130)
         );
  DFF_X1 \REGISTERS_reg[4][56]  ( .D(n6788), .CK(CLK), .Q(n12333), .QN(n16135)
         );
  DFF_X1 \REGISTERS_reg[4][55]  ( .D(n6787), .CK(CLK), .Q(n12334), .QN(n16140)
         );
  DFF_X1 \REGISTERS_reg[4][54]  ( .D(n6786), .CK(CLK), .Q(n12335), .QN(n16145)
         );
  DFF_X1 \REGISTERS_reg[4][53]  ( .D(n6785), .CK(CLK), .Q(n12336), .QN(n16150)
         );
  DFF_X1 \REGISTERS_reg[4][52]  ( .D(n6784), .CK(CLK), .Q(n12337), .QN(n16155)
         );
  DFF_X1 \REGISTERS_reg[4][51]  ( .D(n6783), .CK(CLK), .Q(n12338), .QN(n16160)
         );
  DFF_X1 \REGISTERS_reg[4][50]  ( .D(n6782), .CK(CLK), .Q(n12339), .QN(n16165)
         );
  DFF_X1 \REGISTERS_reg[4][49]  ( .D(n6781), .CK(CLK), .Q(n12340), .QN(n16170)
         );
  DFF_X1 \REGISTERS_reg[4][48]  ( .D(n6780), .CK(CLK), .Q(n12341), .QN(n16175)
         );
  DFF_X1 \REGISTERS_reg[4][47]  ( .D(n6779), .CK(CLK), .Q(n12342), .QN(n16180)
         );
  DFF_X1 \REGISTERS_reg[4][46]  ( .D(n6778), .CK(CLK), .Q(n12343), .QN(n16185)
         );
  DFF_X1 \REGISTERS_reg[4][45]  ( .D(n6777), .CK(CLK), .Q(n12344), .QN(n16190)
         );
  DFF_X1 \REGISTERS_reg[4][44]  ( .D(n6776), .CK(CLK), .Q(n12345), .QN(n16195)
         );
  DFF_X1 \REGISTERS_reg[4][43]  ( .D(n6775), .CK(CLK), .Q(n12346), .QN(n16200)
         );
  DFF_X1 \REGISTERS_reg[4][42]  ( .D(n6774), .CK(CLK), .Q(n12347), .QN(n16205)
         );
  DFF_X1 \REGISTERS_reg[4][41]  ( .D(n6773), .CK(CLK), .Q(n12348), .QN(n16210)
         );
  DFF_X1 \REGISTERS_reg[4][40]  ( .D(n6772), .CK(CLK), .Q(n12349), .QN(n16215)
         );
  DFF_X1 \REGISTERS_reg[4][39]  ( .D(n6771), .CK(CLK), .Q(n12350), .QN(n16220)
         );
  DFF_X1 \REGISTERS_reg[4][38]  ( .D(n6770), .CK(CLK), .Q(n12351), .QN(n16225)
         );
  DFF_X1 \REGISTERS_reg[4][37]  ( .D(n6769), .CK(CLK), .Q(n12352), .QN(n16230)
         );
  DFF_X1 \REGISTERS_reg[4][36]  ( .D(n6768), .CK(CLK), .Q(n12353), .QN(n16235)
         );
  DFF_X1 \REGISTERS_reg[4][35]  ( .D(n6767), .CK(CLK), .Q(n12354), .QN(n16240)
         );
  DFF_X1 \REGISTERS_reg[4][34]  ( .D(n6766), .CK(CLK), .Q(n12355), .QN(n16245)
         );
  DFF_X1 \REGISTERS_reg[4][33]  ( .D(n6765), .CK(CLK), .Q(n12356), .QN(n16250)
         );
  DFF_X1 \REGISTERS_reg[4][32]  ( .D(n6764), .CK(CLK), .Q(n12357), .QN(n16255)
         );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n6763), .CK(CLK), .Q(n12358), .QN(n16260)
         );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n6762), .CK(CLK), .Q(n12359), .QN(n16265)
         );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n6761), .CK(CLK), .Q(n12360), .QN(n16270)
         );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n6760), .CK(CLK), .Q(n12361), .QN(n16275)
         );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n6759), .CK(CLK), .Q(n12362), .QN(n16280)
         );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n6758), .CK(CLK), .Q(n12363), .QN(n16285)
         );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n6757), .CK(CLK), .Q(n12364), .QN(n16290)
         );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n6756), .CK(CLK), .Q(n12365), .QN(n16295)
         );
  DFF_X1 \REGISTERS_reg[1][59]  ( .D(n6983), .CK(CLK), .Q(n12266), .QN(n7877)
         );
  DFF_X1 \REGISTERS_reg[1][58]  ( .D(n6982), .CK(CLK), .Q(n12267), .QN(n7880)
         );
  DFF_X1 \REGISTERS_reg[1][57]  ( .D(n6981), .CK(CLK), .Q(n12268), .QN(n7883)
         );
  DFF_X1 \REGISTERS_reg[1][56]  ( .D(n6980), .CK(CLK), .Q(n12269), .QN(n7886)
         );
  DFF_X1 \REGISTERS_reg[1][55]  ( .D(n6979), .CK(CLK), .Q(n12270), .QN(n7889)
         );
  DFF_X1 \REGISTERS_reg[1][54]  ( .D(n6978), .CK(CLK), .Q(n12271), .QN(n7892)
         );
  DFF_X1 \REGISTERS_reg[1][53]  ( .D(n6977), .CK(CLK), .Q(n12272), .QN(n7895)
         );
  DFF_X1 \REGISTERS_reg[1][52]  ( .D(n6976), .CK(CLK), .Q(n12273), .QN(n7898)
         );
  DFF_X1 \REGISTERS_reg[1][51]  ( .D(n6975), .CK(CLK), .Q(n12274), .QN(n7901)
         );
  DFF_X1 \REGISTERS_reg[1][50]  ( .D(n6974), .CK(CLK), .Q(n12275), .QN(n7904)
         );
  DFF_X1 \REGISTERS_reg[1][49]  ( .D(n6973), .CK(CLK), .Q(n12276), .QN(n7907)
         );
  DFF_X1 \REGISTERS_reg[1][48]  ( .D(n6972), .CK(CLK), .Q(n12277), .QN(n7910)
         );
  DFF_X1 \REGISTERS_reg[1][47]  ( .D(n6971), .CK(CLK), .Q(n12278), .QN(n7913)
         );
  DFF_X1 \REGISTERS_reg[1][46]  ( .D(n6970), .CK(CLK), .Q(n12279), .QN(n7916)
         );
  DFF_X1 \REGISTERS_reg[1][45]  ( .D(n6969), .CK(CLK), .Q(n12280), .QN(n7919)
         );
  DFF_X1 \REGISTERS_reg[1][44]  ( .D(n6968), .CK(CLK), .Q(n12281), .QN(n7922)
         );
  DFF_X1 \REGISTERS_reg[1][43]  ( .D(n6967), .CK(CLK), .Q(n12282), .QN(n7925)
         );
  DFF_X1 \REGISTERS_reg[1][42]  ( .D(n6966), .CK(CLK), .Q(n12283), .QN(n7928)
         );
  DFF_X1 \REGISTERS_reg[1][41]  ( .D(n6965), .CK(CLK), .Q(n12284), .QN(n7931)
         );
  DFF_X1 \REGISTERS_reg[1][40]  ( .D(n6964), .CK(CLK), .Q(n12285), .QN(n7934)
         );
  DFF_X1 \REGISTERS_reg[1][39]  ( .D(n6963), .CK(CLK), .Q(n12286), .QN(n7937)
         );
  DFF_X1 \REGISTERS_reg[1][38]  ( .D(n6962), .CK(CLK), .Q(n12287), .QN(n7940)
         );
  DFF_X1 \REGISTERS_reg[1][37]  ( .D(n6961), .CK(CLK), .Q(n12288), .QN(n7943)
         );
  DFF_X1 \REGISTERS_reg[1][36]  ( .D(n6960), .CK(CLK), .Q(n12289), .QN(n7946)
         );
  DFF_X1 \REGISTERS_reg[1][35]  ( .D(n6959), .CK(CLK), .Q(n12290), .QN(n7949)
         );
  DFF_X1 \REGISTERS_reg[1][34]  ( .D(n6958), .CK(CLK), .Q(n12291), .QN(n7952)
         );
  DFF_X1 \REGISTERS_reg[1][33]  ( .D(n6957), .CK(CLK), .Q(n12292), .QN(n7955)
         );
  DFF_X1 \REGISTERS_reg[1][32]  ( .D(n6956), .CK(CLK), .Q(n12293), .QN(n7958)
         );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n6955), .CK(CLK), .Q(n12294), .QN(n7961)
         );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n6954), .CK(CLK), .Q(n12295), .QN(n7964)
         );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n6953), .CK(CLK), .Q(n12296), .QN(n7967)
         );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n6952), .CK(CLK), .Q(n12297), .QN(n7970)
         );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n6951), .CK(CLK), .Q(n12298), .QN(n7973)
         );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n6950), .CK(CLK), .Q(n12299), .QN(n7976)
         );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n6949), .CK(CLK), .Q(n12300), .QN(n7979)
         );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n6948), .CK(CLK), .Q(n12301), .QN(n7982)
         );
  DFF_X1 \REGISTERS_reg[0][59]  ( .D(n7047), .CK(CLK), .Q(n12202), .QN(n7316)
         );
  DFF_X1 \REGISTERS_reg[0][58]  ( .D(n7046), .CK(CLK), .Q(n12203), .QN(n7318)
         );
  DFF_X1 \REGISTERS_reg[0][57]  ( .D(n7045), .CK(CLK), .Q(n12204), .QN(n7320)
         );
  DFF_X1 \REGISTERS_reg[0][56]  ( .D(n7044), .CK(CLK), .Q(n12205), .QN(n7322)
         );
  DFF_X1 \REGISTERS_reg[0][55]  ( .D(n7043), .CK(CLK), .Q(n12206), .QN(n7324)
         );
  DFF_X1 \REGISTERS_reg[0][54]  ( .D(n7042), .CK(CLK), .Q(n12207), .QN(n7326)
         );
  DFF_X1 \REGISTERS_reg[0][53]  ( .D(n7041), .CK(CLK), .Q(n12208), .QN(n7328)
         );
  DFF_X1 \REGISTERS_reg[0][52]  ( .D(n7040), .CK(CLK), .Q(n12209), .QN(n7330)
         );
  DFF_X1 \REGISTERS_reg[0][51]  ( .D(n7039), .CK(CLK), .Q(n12210), .QN(n7332)
         );
  DFF_X1 \REGISTERS_reg[0][50]  ( .D(n7038), .CK(CLK), .Q(n12211), .QN(n7334)
         );
  DFF_X1 \REGISTERS_reg[0][49]  ( .D(n7037), .CK(CLK), .Q(n12212), .QN(n7336)
         );
  DFF_X1 \REGISTERS_reg[0][48]  ( .D(n7036), .CK(CLK), .Q(n12213), .QN(n7338)
         );
  DFF_X1 \REGISTERS_reg[0][47]  ( .D(n7035), .CK(CLK), .Q(n12214), .QN(n7340)
         );
  DFF_X1 \REGISTERS_reg[0][46]  ( .D(n7034), .CK(CLK), .Q(n12215), .QN(n7342)
         );
  DFF_X1 \REGISTERS_reg[0][45]  ( .D(n7033), .CK(CLK), .Q(n12216), .QN(n7344)
         );
  DFF_X1 \REGISTERS_reg[0][44]  ( .D(n7032), .CK(CLK), .Q(n12217), .QN(n7346)
         );
  DFF_X1 \REGISTERS_reg[0][43]  ( .D(n7031), .CK(CLK), .Q(n12218), .QN(n7348)
         );
  DFF_X1 \REGISTERS_reg[0][42]  ( .D(n7030), .CK(CLK), .Q(n12219), .QN(n7350)
         );
  DFF_X1 \REGISTERS_reg[0][41]  ( .D(n7029), .CK(CLK), .Q(n12220), .QN(n7352)
         );
  DFF_X1 \REGISTERS_reg[0][40]  ( .D(n7028), .CK(CLK), .Q(n12221), .QN(n7354)
         );
  DFF_X1 \REGISTERS_reg[0][39]  ( .D(n7027), .CK(CLK), .Q(n12222), .QN(n7356)
         );
  DFF_X1 \REGISTERS_reg[0][38]  ( .D(n7026), .CK(CLK), .Q(n12223), .QN(n7358)
         );
  DFF_X1 \REGISTERS_reg[0][37]  ( .D(n7025), .CK(CLK), .Q(n12224), .QN(n7360)
         );
  DFF_X1 \REGISTERS_reg[0][36]  ( .D(n7024), .CK(CLK), .Q(n12225), .QN(n7362)
         );
  DFF_X1 \REGISTERS_reg[0][35]  ( .D(n7023), .CK(CLK), .Q(n12226), .QN(n7364)
         );
  DFF_X1 \REGISTERS_reg[0][34]  ( .D(n7022), .CK(CLK), .Q(n12227), .QN(n7366)
         );
  DFF_X1 \REGISTERS_reg[0][33]  ( .D(n7021), .CK(CLK), .Q(n12228), .QN(n7368)
         );
  DFF_X1 \REGISTERS_reg[0][32]  ( .D(n7020), .CK(CLK), .Q(n12229), .QN(n7370)
         );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n7019), .CK(CLK), .Q(n12230), .QN(n7372)
         );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n7018), .CK(CLK), .Q(n12231), .QN(n7374)
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n7017), .CK(CLK), .Q(n12232), .QN(n7376)
         );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n7016), .CK(CLK), .Q(n12233), .QN(n7378)
         );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n7015), .CK(CLK), .Q(n12234), .QN(n7380)
         );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n7014), .CK(CLK), .Q(n12235), .QN(n7382)
         );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n7013), .CK(CLK), .Q(n12236), .QN(n7384)
         );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n7012), .CK(CLK), .Q(n12237), .QN(n7386)
         );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n5219), .CK(CLK), .Q(n13419), .QN(n7689)
         );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n5218), .CK(CLK), .Q(n13420), .QN(n7691)
         );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n5217), .CK(CLK), .Q(n13421), .QN(n7693)
         );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n5216), .CK(CLK), .Q(n13422), .QN(n7695)
         );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n5215), .CK(CLK), .Q(n13423), .QN(n7697)
         );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n5214), .CK(CLK), .Q(n13424), .QN(n7699)
         );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n5213), .CK(CLK), .Q(n13425), .QN(n7701)
         );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n5212), .CK(CLK), .Q(n13426), .QN(n7703)
         );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n5211), .CK(CLK), .Q(n13427), .QN(n7705)
         );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n5210), .CK(CLK), .Q(n13428), .QN(n7707)
         );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n5209), .CK(CLK), .Q(n13429), .QN(n7709)
         );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n5208), .CK(CLK), .Q(n13430), .QN(n7711)
         );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n5207), .CK(CLK), .Q(n13431), .QN(n7713)
         );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n5206), .CK(CLK), .Q(n13432), .QN(n7715)
         );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n5205), .CK(CLK), .Q(n13433), .QN(n7717)
         );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n5204), .CK(CLK), .Q(n13434), .QN(n7719)
         );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n5203), .CK(CLK), .Q(n13435), .QN(n7721)
         );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n5202), .CK(CLK), .Q(n13436), .QN(n7723)
         );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n5201), .CK(CLK), .Q(n13437), .QN(n7725)
         );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n5200), .CK(CLK), .Q(n13438), .QN(n7727)
         );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n5199), .CK(CLK), .Q(n13439), .QN(n7729)
         );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n5198), .CK(CLK), .Q(n13440), .QN(n7731)
         );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n5197), .CK(CLK), .Q(n13441), .QN(n7733)
         );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n5196), .CK(CLK), .Q(n13442), .QN(n7735)
         );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n5411), .CK(CLK), .Q(n13227), .QN(n7284)
         );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n5410), .CK(CLK), .Q(n13228), .QN(n7285)
         );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n5409), .CK(CLK), .Q(n13229), .QN(n7286)
         );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n5408), .CK(CLK), .Q(n13230), .QN(n7287)
         );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n5407), .CK(CLK), .Q(n13231), .QN(n7288)
         );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n5406), .CK(CLK), .Q(n13232), .QN(n7289)
         );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n5405), .CK(CLK), .Q(n13233), .QN(n7290)
         );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n5404), .CK(CLK), .Q(n13234), .QN(n7291)
         );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n5403), .CK(CLK), .Q(n13235), .QN(n7292)
         );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n5402), .CK(CLK), .Q(n13236), .QN(n7293)
         );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n5401), .CK(CLK), .Q(n13237), .QN(n7294)
         );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n5400), .CK(CLK), .Q(n13238), .QN(n7295)
         );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n5399), .CK(CLK), .Q(n13239), .QN(n7296)
         );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n5398), .CK(CLK), .Q(n13240), .QN(n7297)
         );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n5397), .CK(CLK), .Q(n13241), .QN(n7298)
         );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n5396), .CK(CLK), .Q(n13242), .QN(n7299)
         );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n5395), .CK(CLK), .Q(n13243), .QN(n7300)
         );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n5394), .CK(CLK), .Q(n13244), .QN(n7301)
         );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n5393), .CK(CLK), .Q(n13245), .QN(n7302)
         );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n5392), .CK(CLK), .Q(n13246), .QN(n7303)
         );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n5391), .CK(CLK), .Q(n13247), .QN(n7304)
         );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n5390), .CK(CLK), .Q(n13248), .QN(n7305)
         );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n5389), .CK(CLK), .Q(n13249), .QN(n7306)
         );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n5388), .CK(CLK), .Q(n13250), .QN(n7307)
         );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n5475), .CK(CLK), .Q(n13163), .QN(n7987)
         );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n5474), .CK(CLK), .Q(n13164), .QN(n7990)
         );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n5473), .CK(CLK), .Q(n13165), .QN(n7993)
         );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n5472), .CK(CLK), .Q(n13166), .QN(n7996)
         );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n5471), .CK(CLK), .Q(n13167), .QN(n7999)
         );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n5470), .CK(CLK), .Q(n13168), .QN(n8002)
         );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n5469), .CK(CLK), .Q(n13169), .QN(n8005)
         );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n5468), .CK(CLK), .Q(n13170), .QN(n8008)
         );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n5467), .CK(CLK), .Q(n13171), .QN(n8011)
         );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n5466), .CK(CLK), .Q(n13172), .QN(n8014)
         );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n5465), .CK(CLK), .Q(n13173), .QN(n8017)
         );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n5464), .CK(CLK), .Q(n13174), .QN(n8020)
         );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n5463), .CK(CLK), .Q(n13175), .QN(n8023)
         );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n5462), .CK(CLK), .Q(n13176), .QN(n8026)
         );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n5461), .CK(CLK), .Q(n13177), .QN(n8029)
         );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n5460), .CK(CLK), .Q(n13178), .QN(n8032)
         );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n5459), .CK(CLK), .Q(n13179), .QN(n8035)
         );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n5458), .CK(CLK), .Q(n13180), .QN(n8038)
         );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n5457), .CK(CLK), .Q(n13181), .QN(n8041)
         );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n5456), .CK(CLK), .Q(n13182), .QN(n8044)
         );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n5455), .CK(CLK), .Q(n13183), .QN(n8047)
         );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n5454), .CK(CLK), .Q(n13184), .QN(n8050)
         );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n5453), .CK(CLK), .Q(n13185), .QN(n8053)
         );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n5452), .CK(CLK), .Q(n13186), .QN(n8056)
         );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n5603), .CK(CLK), .Q(n13099), .QN(n7389)
         );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n5602), .CK(CLK), .Q(n13100), .QN(n7391)
         );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n5601), .CK(CLK), .Q(n13101), .QN(n7393)
         );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n5600), .CK(CLK), .Q(n13102), .QN(n7395)
         );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n5599), .CK(CLK), .Q(n13103), .QN(n7397)
         );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n5598), .CK(CLK), .Q(n13104), .QN(n7399)
         );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n5597), .CK(CLK), .Q(n13105), .QN(n7401)
         );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n5596), .CK(CLK), .Q(n13106), .QN(n7403)
         );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n5595), .CK(CLK), .Q(n13107), .QN(n7405)
         );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n5594), .CK(CLK), .Q(n13108), .QN(n7407)
         );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n5593), .CK(CLK), .Q(n13109), .QN(n7409)
         );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n5592), .CK(CLK), .Q(n13110), .QN(n7411)
         );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n5591), .CK(CLK), .Q(n13111), .QN(n7413)
         );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n5590), .CK(CLK), .Q(n13112), .QN(n7415)
         );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n5589), .CK(CLK), .Q(n13113), .QN(n7417)
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n5588), .CK(CLK), .Q(n13114), .QN(n7419)
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n5587), .CK(CLK), .Q(n13115), .QN(n7421)
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n5586), .CK(CLK), .Q(n13116), .QN(n7423)
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n5585), .CK(CLK), .Q(n13117), .QN(n7425)
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n5584), .CK(CLK), .Q(n13118), .QN(n7427)
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n5583), .CK(CLK), .Q(n13119), .QN(n7429)
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n5582), .CK(CLK), .Q(n13120), .QN(n7431)
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n5581), .CK(CLK), .Q(n13121), .QN(n7433)
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n5580), .CK(CLK), .Q(n13122), .QN(n7435)
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n6691), .CK(CLK), .Q(n12430), .QN(n7092)
         );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n6690), .CK(CLK), .Q(n12431), .QN(n7093)
         );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n6689), .CK(CLK), .Q(n12432), .QN(n7094)
         );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n6688), .CK(CLK), .Q(n12433), .QN(n7095)
         );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n6687), .CK(CLK), .Q(n12434), .QN(n7096)
         );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n6686), .CK(CLK), .Q(n12435), .QN(n7097)
         );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n6685), .CK(CLK), .Q(n12436), .QN(n7098)
         );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n6684), .CK(CLK), .Q(n12437), .QN(n7099)
         );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n6683), .CK(CLK), .Q(n12438), .QN(n7100)
         );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n6682), .CK(CLK), .Q(n12439), .QN(n7101)
         );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n6681), .CK(CLK), .Q(n12440), .QN(n7102)
         );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n6680), .CK(CLK), .Q(n12441), .QN(n7103)
         );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n6679), .CK(CLK), .Q(n12442), .QN(n7104)
         );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n6678), .CK(CLK), .Q(n12443), .QN(n7105)
         );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n6677), .CK(CLK), .Q(n12444), .QN(n7106)
         );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n6676), .CK(CLK), .Q(n12445), .QN(n7107)
         );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n6675), .CK(CLK), .Q(n12446), .QN(n7108)
         );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n6674), .CK(CLK), .Q(n12447), .QN(n7109)
         );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n6673), .CK(CLK), .Q(n12448), .QN(n7110)
         );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n6672), .CK(CLK), .Q(n12449), .QN(n7111)
         );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n6671), .CK(CLK), .Q(n12450), .QN(n7112)
         );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n6670), .CK(CLK), .Q(n12451), .QN(n7113)
         );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n6669), .CK(CLK), .Q(n12452), .QN(n7114)
         );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n6668), .CK(CLK), .Q(n12453), .QN(n7115)
         );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n6755), .CK(CLK), .Q(n12366), .QN(n16300)
         );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n6754), .CK(CLK), .Q(n12367), .QN(n16305)
         );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n6753), .CK(CLK), .Q(n12368), .QN(n16310)
         );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n6752), .CK(CLK), .Q(n12369), .QN(n16315)
         );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n6751), .CK(CLK), .Q(n12370), .QN(n16320)
         );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n6750), .CK(CLK), .Q(n12371), .QN(n16325)
         );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n6749), .CK(CLK), .Q(n12372), .QN(n16330)
         );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n6748), .CK(CLK), .Q(n12373), .QN(n16335)
         );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n6747), .CK(CLK), .Q(n12374), .QN(n16340)
         );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n6746), .CK(CLK), .Q(n12375), .QN(n16345)
         );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n6745), .CK(CLK), .Q(n12376), .QN(n16350)
         );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n6744), .CK(CLK), .Q(n12377), .QN(n16355)
         );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n6743), .CK(CLK), .Q(n12378), .QN(n16360)
         );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n6742), .CK(CLK), .Q(n12379), .QN(n16365)
         );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n6741), .CK(CLK), .Q(n12380), .QN(n16370)
         );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n6740), .CK(CLK), .Q(n12381), .QN(n16375)
         );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n6739), .CK(CLK), .Q(n12382), .QN(n16380)
         );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n6738), .CK(CLK), .Q(n12383), .QN(n16385)
         );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n6737), .CK(CLK), .Q(n12384), .QN(n16390)
         );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n6736), .CK(CLK), .Q(n12385), .QN(n16395)
         );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n6735), .CK(CLK), .Q(n12386), .QN(n16400)
         );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n6734), .CK(CLK), .Q(n12387), .QN(n16405)
         );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n6733), .CK(CLK), .Q(n12388), .QN(n16410)
         );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n6732), .CK(CLK), .Q(n12389), .QN(n16415)
         );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n6947), .CK(CLK), .Q(n12302), .QN(n7985)
         );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n6946), .CK(CLK), .Q(n12303), .QN(n7988)
         );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n6945), .CK(CLK), .Q(n12304), .QN(n7991)
         );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n6944), .CK(CLK), .Q(n12305), .QN(n7994)
         );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n6943), .CK(CLK), .Q(n12306), .QN(n7997)
         );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n6942), .CK(CLK), .Q(n12307), .QN(n8000)
         );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n6941), .CK(CLK), .Q(n12308), .QN(n8003)
         );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n6940), .CK(CLK), .Q(n12309), .QN(n8006)
         );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n6939), .CK(CLK), .Q(n12310), .QN(n8009)
         );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n6938), .CK(CLK), .Q(n12311), .QN(n8012)
         );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n6937), .CK(CLK), .Q(n12312), .QN(n8015)
         );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n6936), .CK(CLK), .Q(n12313), .QN(n8018)
         );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n6935), .CK(CLK), .Q(n12314), .QN(n8021)
         );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n6934), .CK(CLK), .Q(n12315), .QN(n8024)
         );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n6933), .CK(CLK), .Q(n12316), .QN(n8027)
         );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n6932), .CK(CLK), .Q(n12317), .QN(n8030)
         );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n6931), .CK(CLK), .Q(n12318), .QN(n8033)
         );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n6930), .CK(CLK), .Q(n12319), .QN(n8036)
         );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n6929), .CK(CLK), .Q(n12320), .QN(n8039)
         );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n6928), .CK(CLK), .Q(n12321), .QN(n8042)
         );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n6927), .CK(CLK), .Q(n12322), .QN(n8045)
         );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n6926), .CK(CLK), .Q(n12323), .QN(n8048)
         );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n6925), .CK(CLK), .Q(n12324), .QN(n8051)
         );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n6924), .CK(CLK), .Q(n12325), .QN(n8054)
         );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n7011), .CK(CLK), .Q(n12238), .QN(n7388)
         );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n7010), .CK(CLK), .Q(n12239), .QN(n7390)
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n7009), .CK(CLK), .Q(n12240), .QN(n7392)
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n7008), .CK(CLK), .Q(n12241), .QN(n7394)
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n7007), .CK(CLK), .Q(n12242), .QN(n7396)
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n7006), .CK(CLK), .Q(n12243), .QN(n7398)
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n7005), .CK(CLK), .Q(n12244), .QN(n7400)
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n7004), .CK(CLK), .Q(n12245), .QN(n7402)
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n7003), .CK(CLK), .Q(n12246), .QN(n7404)
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n7002), .CK(CLK), .Q(n12247), .QN(n7406)
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n7001), .CK(CLK), .Q(n12248), .QN(n7408)
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n7000), .CK(CLK), .Q(n12249), .QN(n7410)
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n6999), .CK(CLK), .Q(n12250), .QN(n7412)
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n6998), .CK(CLK), .Q(n12251), .QN(n7414)
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n6997), .CK(CLK), .Q(n12252), .QN(n7416)
         );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n6996), .CK(CLK), .Q(n12253), .QN(n7418)
         );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n6995), .CK(CLK), .Q(n12254), .QN(n7420)
         );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n6994), .CK(CLK), .Q(n12255), .QN(n7422)
         );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n6993), .CK(CLK), .Q(n12256), .QN(n7424)
         );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n6992), .CK(CLK), .Q(n12257), .QN(n7426)
         );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n6991), .CK(CLK), .Q(n12258), .QN(n7428)
         );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n6990), .CK(CLK), .Q(n12259), .QN(n7430)
         );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n6989), .CK(CLK), .Q(n12260), .QN(n7432)
         );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n6988), .CK(CLK), .Q(n12261), .QN(n7434)
         );
  DFF_X1 \REGISTERS_reg[29][63]  ( .D(n5195), .CK(CLK), .QN(n7737) );
  DFF_X1 \REGISTERS_reg[12][63]  ( .D(n6283), .CK(CLK), .QN(n12710) );
  DFF_X1 \REGISTERS_reg[12][62]  ( .D(n6282), .CK(CLK), .QN(n12711) );
  DFF_X1 \REGISTERS_reg[12][61]  ( .D(n6281), .CK(CLK), .QN(n12712) );
  DFF_X1 \REGISTERS_reg[12][60]  ( .D(n6280), .CK(CLK), .QN(n12713) );
  DFF_X1 \REGISTERS_reg[10][63]  ( .D(n6411), .CK(CLK), .QN(n12582) );
  DFF_X1 \REGISTERS_reg[10][62]  ( .D(n6410), .CK(CLK), .QN(n12583) );
  DFF_X1 \REGISTERS_reg[10][61]  ( .D(n6409), .CK(CLK), .QN(n12584) );
  DFF_X1 \REGISTERS_reg[10][60]  ( .D(n6408), .CK(CLK), .QN(n12585) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n6029), .CK(CLK), .QN(n12801) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n6028), .CK(CLK), .QN(n12802) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n6056), .CK(CLK), .QN(n12774) );
  DFF_X1 \REGISTERS_reg[12][59]  ( .D(n6279), .CK(CLK), .QN(n12714) );
  DFF_X1 \REGISTERS_reg[12][58]  ( .D(n6278), .CK(CLK), .QN(n12715) );
  DFF_X1 \REGISTERS_reg[12][57]  ( .D(n6277), .CK(CLK), .QN(n12716) );
  DFF_X1 \REGISTERS_reg[12][56]  ( .D(n6276), .CK(CLK), .QN(n12717) );
  DFF_X1 \REGISTERS_reg[12][55]  ( .D(n6275), .CK(CLK), .QN(n12718) );
  DFF_X1 \REGISTERS_reg[12][54]  ( .D(n6274), .CK(CLK), .QN(n12719) );
  DFF_X1 \REGISTERS_reg[12][53]  ( .D(n6273), .CK(CLK), .QN(n12720) );
  DFF_X1 \REGISTERS_reg[12][52]  ( .D(n6272), .CK(CLK), .QN(n12721) );
  DFF_X1 \REGISTERS_reg[12][51]  ( .D(n6271), .CK(CLK), .QN(n12722) );
  DFF_X1 \REGISTERS_reg[12][50]  ( .D(n6270), .CK(CLK), .QN(n12723) );
  DFF_X1 \REGISTERS_reg[12][49]  ( .D(n6269), .CK(CLK), .QN(n12724) );
  DFF_X1 \REGISTERS_reg[12][48]  ( .D(n6268), .CK(CLK), .QN(n12725) );
  DFF_X1 \REGISTERS_reg[12][47]  ( .D(n6267), .CK(CLK), .QN(n12726) );
  DFF_X1 \REGISTERS_reg[12][46]  ( .D(n6266), .CK(CLK), .QN(n12727) );
  DFF_X1 \REGISTERS_reg[12][45]  ( .D(n6265), .CK(CLK), .QN(n12728) );
  DFF_X1 \REGISTERS_reg[12][44]  ( .D(n6264), .CK(CLK), .QN(n12729) );
  DFF_X1 \REGISTERS_reg[12][43]  ( .D(n6263), .CK(CLK), .QN(n12730) );
  DFF_X1 \REGISTERS_reg[12][42]  ( .D(n6262), .CK(CLK), .QN(n12731) );
  DFF_X1 \REGISTERS_reg[12][41]  ( .D(n6261), .CK(CLK), .QN(n12732) );
  DFF_X1 \REGISTERS_reg[12][40]  ( .D(n6260), .CK(CLK), .QN(n12733) );
  DFF_X1 \REGISTERS_reg[12][39]  ( .D(n6259), .CK(CLK), .QN(n12734) );
  DFF_X1 \REGISTERS_reg[12][38]  ( .D(n6258), .CK(CLK), .QN(n12735) );
  DFF_X1 \REGISTERS_reg[12][37]  ( .D(n6257), .CK(CLK), .QN(n12736) );
  DFF_X1 \REGISTERS_reg[12][36]  ( .D(n6256), .CK(CLK), .QN(n12737) );
  DFF_X1 \REGISTERS_reg[12][35]  ( .D(n6255), .CK(CLK), .QN(n12738) );
  DFF_X1 \REGISTERS_reg[12][34]  ( .D(n6254), .CK(CLK), .QN(n12739) );
  DFF_X1 \REGISTERS_reg[12][33]  ( .D(n6253), .CK(CLK), .QN(n12740) );
  DFF_X1 \REGISTERS_reg[12][32]  ( .D(n6252), .CK(CLK), .QN(n12741) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n6251), .CK(CLK), .QN(n12742) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n6250), .CK(CLK), .QN(n12743) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n6249), .CK(CLK), .QN(n12744) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n6248), .CK(CLK), .QN(n12745) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n6247), .CK(CLK), .QN(n12746) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n6246), .CK(CLK), .QN(n12747) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n6245), .CK(CLK), .QN(n12748) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n6244), .CK(CLK), .QN(n12749) );
  DFF_X1 \REGISTERS_reg[10][59]  ( .D(n6407), .CK(CLK), .QN(n12586) );
  DFF_X1 \REGISTERS_reg[10][58]  ( .D(n6406), .CK(CLK), .QN(n12587) );
  DFF_X1 \REGISTERS_reg[10][57]  ( .D(n6405), .CK(CLK), .QN(n12588) );
  DFF_X1 \REGISTERS_reg[10][56]  ( .D(n6404), .CK(CLK), .QN(n12589) );
  DFF_X1 \REGISTERS_reg[10][55]  ( .D(n6403), .CK(CLK), .QN(n12590) );
  DFF_X1 \REGISTERS_reg[10][54]  ( .D(n6402), .CK(CLK), .QN(n12591) );
  DFF_X1 \REGISTERS_reg[10][53]  ( .D(n6401), .CK(CLK), .QN(n12592) );
  DFF_X1 \REGISTERS_reg[10][52]  ( .D(n6400), .CK(CLK), .QN(n12593) );
  DFF_X1 \REGISTERS_reg[10][51]  ( .D(n6399), .CK(CLK), .QN(n12594) );
  DFF_X1 \REGISTERS_reg[10][50]  ( .D(n6398), .CK(CLK), .QN(n12595) );
  DFF_X1 \REGISTERS_reg[10][49]  ( .D(n6397), .CK(CLK), .QN(n12596) );
  DFF_X1 \REGISTERS_reg[10][48]  ( .D(n6396), .CK(CLK), .QN(n12597) );
  DFF_X1 \REGISTERS_reg[10][47]  ( .D(n6395), .CK(CLK), .QN(n12598) );
  DFF_X1 \REGISTERS_reg[10][46]  ( .D(n6394), .CK(CLK), .QN(n12599) );
  DFF_X1 \REGISTERS_reg[10][45]  ( .D(n6393), .CK(CLK), .QN(n12600) );
  DFF_X1 \REGISTERS_reg[10][44]  ( .D(n6392), .CK(CLK), .QN(n12601) );
  DFF_X1 \REGISTERS_reg[10][43]  ( .D(n6391), .CK(CLK), .QN(n12602) );
  DFF_X1 \REGISTERS_reg[10][42]  ( .D(n6390), .CK(CLK), .QN(n12603) );
  DFF_X1 \REGISTERS_reg[10][41]  ( .D(n6389), .CK(CLK), .QN(n12604) );
  DFF_X1 \REGISTERS_reg[10][40]  ( .D(n6388), .CK(CLK), .QN(n12605) );
  DFF_X1 \REGISTERS_reg[10][39]  ( .D(n6387), .CK(CLK), .QN(n12606) );
  DFF_X1 \REGISTERS_reg[10][38]  ( .D(n6386), .CK(CLK), .QN(n12607) );
  DFF_X1 \REGISTERS_reg[10][37]  ( .D(n6385), .CK(CLK), .QN(n12608) );
  DFF_X1 \REGISTERS_reg[10][36]  ( .D(n6384), .CK(CLK), .QN(n12609) );
  DFF_X1 \REGISTERS_reg[10][35]  ( .D(n6383), .CK(CLK), .QN(n12610) );
  DFF_X1 \REGISTERS_reg[10][34]  ( .D(n6382), .CK(CLK), .QN(n12611) );
  DFF_X1 \REGISTERS_reg[10][33]  ( .D(n6381), .CK(CLK), .QN(n12612) );
  DFF_X1 \REGISTERS_reg[10][32]  ( .D(n6380), .CK(CLK), .QN(n12613) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n6379), .CK(CLK), .QN(n12614) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n6378), .CK(CLK), .QN(n12615) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n6377), .CK(CLK), .QN(n12616) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n6376), .CK(CLK), .QN(n12617) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n6375), .CK(CLK), .QN(n12618) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n6374), .CK(CLK), .QN(n12619) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n6373), .CK(CLK), .QN(n12620) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n6372), .CK(CLK), .QN(n12621) );
  DFF_X1 \REGISTERS_reg[31][63]  ( .D(n5067), .CK(CLK), .QN(n13507) );
  DFF_X1 \REGISTERS_reg[31][62]  ( .D(n5066), .CK(CLK), .QN(n13508) );
  DFF_X1 \REGISTERS_reg[31][61]  ( .D(n5065), .CK(CLK), .QN(n13509) );
  DFF_X1 \REGISTERS_reg[31][60]  ( .D(n5064), .CK(CLK), .QN(n13510) );
  DFF_X1 \REGISTERS_reg[30][63]  ( .D(n5131), .CK(CLK), .QN(n13443) );
  DFF_X1 \REGISTERS_reg[30][62]  ( .D(n5130), .CK(CLK), .QN(n13444) );
  DFF_X1 \REGISTERS_reg[30][61]  ( .D(n5129), .CK(CLK), .QN(n13445) );
  DFF_X1 \REGISTERS_reg[30][60]  ( .D(n5128), .CK(CLK), .QN(n13446) );
  DFF_X1 \REGISTERS_reg[21][63]  ( .D(n5707), .CK(CLK), .QN(n12995) );
  DFF_X1 \REGISTERS_reg[21][62]  ( .D(n5706), .CK(CLK), .QN(n12996) );
  DFF_X1 \REGISTERS_reg[21][61]  ( .D(n5705), .CK(CLK), .QN(n12997) );
  DFF_X1 \REGISTERS_reg[21][60]  ( .D(n5704), .CK(CLK), .QN(n12998) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n6243), .CK(CLK), .QN(n12750) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n6242), .CK(CLK), .QN(n12751) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n6241), .CK(CLK), .QN(n12752) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n6240), .CK(CLK), .QN(n12753) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n6239), .CK(CLK), .QN(n12754) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n6238), .CK(CLK), .QN(n12755) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n6237), .CK(CLK), .QN(n12756) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n6236), .CK(CLK), .QN(n12757) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n6235), .CK(CLK), .QN(n12758) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n6234), .CK(CLK), .QN(n12759) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n6233), .CK(CLK), .QN(n12760) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n6232), .CK(CLK), .QN(n12761) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n6231), .CK(CLK), .QN(n12762) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n6230), .CK(CLK), .QN(n12763) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n6229), .CK(CLK), .QN(n12764) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n6228), .CK(CLK), .QN(n12765) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n6227), .CK(CLK), .QN(n12766) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n6226), .CK(CLK), .QN(n12767) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n6225), .CK(CLK), .QN(n12768) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n6224), .CK(CLK), .QN(n12769) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n6223), .CK(CLK), .QN(n12770) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n6222), .CK(CLK), .QN(n12771) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n6221), .CK(CLK), .QN(n12772) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n6220), .CK(CLK), .QN(n12773) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n6371), .CK(CLK), .QN(n12622) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n6370), .CK(CLK), .QN(n12623) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n6369), .CK(CLK), .QN(n12624) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n6368), .CK(CLK), .QN(n12625) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n6367), .CK(CLK), .QN(n12626) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n6366), .CK(CLK), .QN(n12627) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n6365), .CK(CLK), .QN(n12628) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n6364), .CK(CLK), .QN(n12629) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n6363), .CK(CLK), .QN(n12630) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n6362), .CK(CLK), .QN(n12631) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n6361), .CK(CLK), .QN(n12632) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n6360), .CK(CLK), .QN(n12633) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n6359), .CK(CLK), .QN(n12634) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n6358), .CK(CLK), .QN(n12635) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n6357), .CK(CLK), .QN(n12636) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n6356), .CK(CLK), .QN(n12637) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n6355), .CK(CLK), .QN(n12638) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n6354), .CK(CLK), .QN(n12639) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n6353), .CK(CLK), .QN(n12640) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n6352), .CK(CLK), .QN(n12641) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n6351), .CK(CLK), .QN(n12642) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n6350), .CK(CLK), .QN(n12643) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n6349), .CK(CLK), .QN(n12644) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n6348), .CK(CLK), .QN(n12645) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n6055), .CK(CLK), .QN(n12775) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n6054), .CK(CLK), .QN(n12776) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n6053), .CK(CLK), .QN(n12777) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n6052), .CK(CLK), .QN(n12778) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n6051), .CK(CLK), .QN(n12779) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n6050), .CK(CLK), .QN(n12780) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n6049), .CK(CLK), .QN(n12781) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n6048), .CK(CLK), .QN(n12782) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n6047), .CK(CLK), .QN(n12783) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n6046), .CK(CLK), .QN(n12784) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n6045), .CK(CLK), .QN(n12785) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n6044), .CK(CLK), .QN(n12786) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n6043), .CK(CLK), .QN(n12787) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n6042), .CK(CLK), .QN(n12788) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n6041), .CK(CLK), .QN(n12789) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n6040), .CK(CLK), .QN(n12790) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n6039), .CK(CLK), .QN(n12791) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n6038), .CK(CLK), .QN(n12792) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n6037), .CK(CLK), .QN(n12793) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n6036), .CK(CLK), .QN(n12794) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n6035), .CK(CLK), .QN(n12795) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n6034), .CK(CLK), .QN(n12796) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n6033), .CK(CLK), .QN(n12797) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n6032), .CK(CLK), .QN(n12798) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n6031), .CK(CLK), .QN(n12799) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n6030), .CK(CLK), .QN(n12800) );
  DFF_X1 \REGISTERS_reg[31][59]  ( .D(n5063), .CK(CLK), .QN(n13511) );
  DFF_X1 \REGISTERS_reg[31][58]  ( .D(n5062), .CK(CLK), .QN(n13512) );
  DFF_X1 \REGISTERS_reg[31][57]  ( .D(n5061), .CK(CLK), .QN(n13513) );
  DFF_X1 \REGISTERS_reg[31][56]  ( .D(n5060), .CK(CLK), .QN(n13514) );
  DFF_X1 \REGISTERS_reg[31][55]  ( .D(n5059), .CK(CLK), .QN(n13515) );
  DFF_X1 \REGISTERS_reg[31][54]  ( .D(n5058), .CK(CLK), .QN(n13516) );
  DFF_X1 \REGISTERS_reg[31][53]  ( .D(n5057), .CK(CLK), .QN(n13517) );
  DFF_X1 \REGISTERS_reg[31][52]  ( .D(n5056), .CK(CLK), .QN(n13518) );
  DFF_X1 \REGISTERS_reg[31][51]  ( .D(n5055), .CK(CLK), .QN(n13519) );
  DFF_X1 \REGISTERS_reg[31][50]  ( .D(n5054), .CK(CLK), .QN(n13520) );
  DFF_X1 \REGISTERS_reg[31][49]  ( .D(n5053), .CK(CLK), .QN(n13521) );
  DFF_X1 \REGISTERS_reg[31][48]  ( .D(n5052), .CK(CLK), .QN(n13522) );
  DFF_X1 \REGISTERS_reg[31][47]  ( .D(n5051), .CK(CLK), .QN(n13523) );
  DFF_X1 \REGISTERS_reg[31][46]  ( .D(n5050), .CK(CLK), .QN(n13524) );
  DFF_X1 \REGISTERS_reg[31][45]  ( .D(n5049), .CK(CLK), .QN(n13525) );
  DFF_X1 \REGISTERS_reg[31][44]  ( .D(n5048), .CK(CLK), .QN(n13526) );
  DFF_X1 \REGISTERS_reg[31][43]  ( .D(n5047), .CK(CLK), .QN(n13527) );
  DFF_X1 \REGISTERS_reg[31][42]  ( .D(n5046), .CK(CLK), .QN(n13528) );
  DFF_X1 \REGISTERS_reg[31][41]  ( .D(n5045), .CK(CLK), .QN(n13529) );
  DFF_X1 \REGISTERS_reg[31][40]  ( .D(n5044), .CK(CLK), .QN(n13530) );
  DFF_X1 \REGISTERS_reg[31][39]  ( .D(n5043), .CK(CLK), .QN(n13531) );
  DFF_X1 \REGISTERS_reg[31][38]  ( .D(n5042), .CK(CLK), .QN(n13532) );
  DFF_X1 \REGISTERS_reg[31][37]  ( .D(n5041), .CK(CLK), .QN(n13533) );
  DFF_X1 \REGISTERS_reg[31][36]  ( .D(n5040), .CK(CLK), .QN(n13534) );
  DFF_X1 \REGISTERS_reg[31][35]  ( .D(n5039), .CK(CLK), .QN(n13535) );
  DFF_X1 \REGISTERS_reg[31][34]  ( .D(n5038), .CK(CLK), .QN(n13536) );
  DFF_X1 \REGISTERS_reg[31][33]  ( .D(n5037), .CK(CLK), .QN(n13537) );
  DFF_X1 \REGISTERS_reg[31][32]  ( .D(n5036), .CK(CLK), .QN(n13538) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n5035), .CK(CLK), .QN(n13539) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n5034), .CK(CLK), .QN(n13540) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n5033), .CK(CLK), .QN(n13541) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n5032), .CK(CLK), .QN(n13542) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n5031), .CK(CLK), .QN(n13543) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n5030), .CK(CLK), .QN(n13544) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n5029), .CK(CLK), .QN(n13545) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n5028), .CK(CLK), .QN(n13546) );
  DFF_X1 \REGISTERS_reg[30][59]  ( .D(n5127), .CK(CLK), .QN(n13447) );
  DFF_X1 \REGISTERS_reg[30][58]  ( .D(n5126), .CK(CLK), .QN(n13448) );
  DFF_X1 \REGISTERS_reg[30][57]  ( .D(n5125), .CK(CLK), .QN(n13449) );
  DFF_X1 \REGISTERS_reg[30][56]  ( .D(n5124), .CK(CLK), .QN(n13450) );
  DFF_X1 \REGISTERS_reg[30][55]  ( .D(n5123), .CK(CLK), .QN(n13451) );
  DFF_X1 \REGISTERS_reg[30][54]  ( .D(n5122), .CK(CLK), .QN(n13452) );
  DFF_X1 \REGISTERS_reg[30][53]  ( .D(n5121), .CK(CLK), .QN(n13453) );
  DFF_X1 \REGISTERS_reg[30][52]  ( .D(n5120), .CK(CLK), .QN(n13454) );
  DFF_X1 \REGISTERS_reg[30][51]  ( .D(n5119), .CK(CLK), .QN(n13455) );
  DFF_X1 \REGISTERS_reg[30][50]  ( .D(n5118), .CK(CLK), .QN(n13456) );
  DFF_X1 \REGISTERS_reg[30][49]  ( .D(n5117), .CK(CLK), .QN(n13457) );
  DFF_X1 \REGISTERS_reg[30][48]  ( .D(n5116), .CK(CLK), .QN(n13458) );
  DFF_X1 \REGISTERS_reg[30][47]  ( .D(n5115), .CK(CLK), .QN(n13459) );
  DFF_X1 \REGISTERS_reg[30][46]  ( .D(n5114), .CK(CLK), .QN(n13460) );
  DFF_X1 \REGISTERS_reg[30][45]  ( .D(n5113), .CK(CLK), .QN(n13461) );
  DFF_X1 \REGISTERS_reg[30][44]  ( .D(n5112), .CK(CLK), .QN(n13462) );
  DFF_X1 \REGISTERS_reg[30][43]  ( .D(n5111), .CK(CLK), .QN(n13463) );
  DFF_X1 \REGISTERS_reg[30][42]  ( .D(n5110), .CK(CLK), .QN(n13464) );
  DFF_X1 \REGISTERS_reg[30][41]  ( .D(n5109), .CK(CLK), .QN(n13465) );
  DFF_X1 \REGISTERS_reg[30][40]  ( .D(n5108), .CK(CLK), .QN(n13466) );
  DFF_X1 \REGISTERS_reg[30][39]  ( .D(n5107), .CK(CLK), .QN(n13467) );
  DFF_X1 \REGISTERS_reg[30][38]  ( .D(n5106), .CK(CLK), .QN(n13468) );
  DFF_X1 \REGISTERS_reg[30][37]  ( .D(n5105), .CK(CLK), .QN(n13469) );
  DFF_X1 \REGISTERS_reg[30][36]  ( .D(n5104), .CK(CLK), .QN(n13470) );
  DFF_X1 \REGISTERS_reg[30][35]  ( .D(n5103), .CK(CLK), .QN(n13471) );
  DFF_X1 \REGISTERS_reg[30][34]  ( .D(n5102), .CK(CLK), .QN(n13472) );
  DFF_X1 \REGISTERS_reg[30][33]  ( .D(n5101), .CK(CLK), .QN(n13473) );
  DFF_X1 \REGISTERS_reg[30][32]  ( .D(n5100), .CK(CLK), .QN(n13474) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n5099), .CK(CLK), .QN(n13475) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n5098), .CK(CLK), .QN(n13476) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n5097), .CK(CLK), .QN(n13477) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n5096), .CK(CLK), .QN(n13478) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n5095), .CK(CLK), .QN(n13479) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n5094), .CK(CLK), .QN(n13480) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n5093), .CK(CLK), .QN(n13481) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n5092), .CK(CLK), .QN(n13482) );
  DFF_X1 \REGISTERS_reg[21][59]  ( .D(n5703), .CK(CLK), .QN(n12999) );
  DFF_X1 \REGISTERS_reg[21][58]  ( .D(n5702), .CK(CLK), .QN(n13000) );
  DFF_X1 \REGISTERS_reg[21][57]  ( .D(n5701), .CK(CLK), .QN(n13001) );
  DFF_X1 \REGISTERS_reg[21][56]  ( .D(n5700), .CK(CLK), .QN(n13002) );
  DFF_X1 \REGISTERS_reg[21][55]  ( .D(n5699), .CK(CLK), .QN(n13003) );
  DFF_X1 \REGISTERS_reg[21][54]  ( .D(n5698), .CK(CLK), .QN(n13004) );
  DFF_X1 \REGISTERS_reg[21][53]  ( .D(n5697), .CK(CLK), .QN(n13005) );
  DFF_X1 \REGISTERS_reg[21][52]  ( .D(n5696), .CK(CLK), .QN(n13006) );
  DFF_X1 \REGISTERS_reg[21][51]  ( .D(n5695), .CK(CLK), .QN(n13007) );
  DFF_X1 \REGISTERS_reg[21][50]  ( .D(n5694), .CK(CLK), .QN(n13008) );
  DFF_X1 \REGISTERS_reg[21][49]  ( .D(n5693), .CK(CLK), .QN(n13009) );
  DFF_X1 \REGISTERS_reg[21][48]  ( .D(n5692), .CK(CLK), .QN(n13010) );
  DFF_X1 \REGISTERS_reg[21][47]  ( .D(n5691), .CK(CLK), .QN(n13011) );
  DFF_X1 \REGISTERS_reg[21][46]  ( .D(n5690), .CK(CLK), .QN(n13012) );
  DFF_X1 \REGISTERS_reg[21][45]  ( .D(n5689), .CK(CLK), .QN(n13013) );
  DFF_X1 \REGISTERS_reg[21][44]  ( .D(n5688), .CK(CLK), .QN(n13014) );
  DFF_X1 \REGISTERS_reg[21][43]  ( .D(n5687), .CK(CLK), .QN(n13015) );
  DFF_X1 \REGISTERS_reg[21][42]  ( .D(n5686), .CK(CLK), .QN(n13016) );
  DFF_X1 \REGISTERS_reg[21][41]  ( .D(n5685), .CK(CLK), .QN(n13017) );
  DFF_X1 \REGISTERS_reg[21][40]  ( .D(n5684), .CK(CLK), .QN(n13018) );
  DFF_X1 \REGISTERS_reg[21][39]  ( .D(n5683), .CK(CLK), .QN(n13019) );
  DFF_X1 \REGISTERS_reg[21][38]  ( .D(n5682), .CK(CLK), .QN(n13020) );
  DFF_X1 \REGISTERS_reg[21][37]  ( .D(n5681), .CK(CLK), .QN(n13021) );
  DFF_X1 \REGISTERS_reg[21][36]  ( .D(n5680), .CK(CLK), .QN(n13022) );
  DFF_X1 \REGISTERS_reg[21][35]  ( .D(n5679), .CK(CLK), .QN(n13023) );
  DFF_X1 \REGISTERS_reg[21][34]  ( .D(n5678), .CK(CLK), .QN(n13024) );
  DFF_X1 \REGISTERS_reg[21][33]  ( .D(n5677), .CK(CLK), .QN(n13025) );
  DFF_X1 \REGISTERS_reg[21][32]  ( .D(n5676), .CK(CLK), .QN(n13026) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n5675), .CK(CLK), .QN(n13027) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n5674), .CK(CLK), .QN(n13028) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n5673), .CK(CLK), .QN(n13029) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n5672), .CK(CLK), .QN(n13030) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n5671), .CK(CLK), .QN(n13031) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n5670), .CK(CLK), .QN(n13032) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n5669), .CK(CLK), .QN(n13033) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n5668), .CK(CLK), .QN(n13034) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n5027), .CK(CLK), .QN(n13547) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n5026), .CK(CLK), .QN(n13548) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n5025), .CK(CLK), .QN(n13549) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n5024), .CK(CLK), .QN(n13550) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n5023), .CK(CLK), .QN(n13551) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n5022), .CK(CLK), .QN(n13552) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n5021), .CK(CLK), .QN(n13553) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n5020), .CK(CLK), .QN(n13554) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n5019), .CK(CLK), .QN(n13555) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n5018), .CK(CLK), .QN(n13556) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n5017), .CK(CLK), .QN(n13557) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n5016), .CK(CLK), .QN(n13558) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n5015), .CK(CLK), .QN(n13559) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n5014), .CK(CLK), .QN(n13560) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n5013), .CK(CLK), .QN(n13561) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n5012), .CK(CLK), .QN(n13562) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n5011), .CK(CLK), .QN(n13563) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n5010), .CK(CLK), .QN(n13564) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n5009), .CK(CLK), .QN(n13565) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n5008), .CK(CLK), .QN(n13566) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n5007), .CK(CLK), .QN(n13567) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n5006), .CK(CLK), .QN(n13568) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n5005), .CK(CLK), .QN(n13569) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n5004), .CK(CLK), .QN(n13570) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n5091), .CK(CLK), .QN(n13483) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n5090), .CK(CLK), .QN(n13484) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n5089), .CK(CLK), .QN(n13485) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n5088), .CK(CLK), .QN(n13486) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n5087), .CK(CLK), .QN(n13487) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n5086), .CK(CLK), .QN(n13488) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n5085), .CK(CLK), .QN(n13489) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n5084), .CK(CLK), .QN(n13490) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n5083), .CK(CLK), .QN(n13491) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n5082), .CK(CLK), .QN(n13492) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n5081), .CK(CLK), .QN(n13493) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n5080), .CK(CLK), .QN(n13494) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n5079), .CK(CLK), .QN(n13495) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n5078), .CK(CLK), .QN(n13496) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n5077), .CK(CLK), .QN(n13497) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n5076), .CK(CLK), .QN(n13498) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n5075), .CK(CLK), .QN(n13499) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n5074), .CK(CLK), .QN(n13500) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n5073), .CK(CLK), .QN(n13501) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n5072), .CK(CLK), .QN(n13502) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n5071), .CK(CLK), .QN(n13503) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n5070), .CK(CLK), .QN(n13504) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n5069), .CK(CLK), .QN(n13505) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n5068), .CK(CLK), .QN(n13506) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n5667), .CK(CLK), .QN(n13035) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n5666), .CK(CLK), .QN(n13036) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n5665), .CK(CLK), .QN(n13037) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n5664), .CK(CLK), .QN(n13038) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n5663), .CK(CLK), .QN(n13039) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n5662), .CK(CLK), .QN(n13040) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n5661), .CK(CLK), .QN(n13041) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n5660), .CK(CLK), .QN(n13042) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n5659), .CK(CLK), .QN(n13043) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n5658), .CK(CLK), .QN(n13044) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n5657), .CK(CLK), .QN(n13045) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n5656), .CK(CLK), .QN(n13046) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n5655), .CK(CLK), .QN(n13047) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n5654), .CK(CLK), .QN(n13048) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n5653), .CK(CLK), .QN(n13049) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n5652), .CK(CLK), .QN(n13050) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n5651), .CK(CLK), .QN(n13051) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n5650), .CK(CLK), .QN(n13052) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n5649), .CK(CLK), .QN(n13053) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n5648), .CK(CLK), .QN(n13054) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n5647), .CK(CLK), .QN(n13055) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n5646), .CK(CLK), .QN(n13056) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n5645), .CK(CLK), .QN(n13057) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n5644), .CK(CLK), .QN(n13058) );
  DFF_X1 \REGISTERS_reg[9][63]  ( .D(n6475), .CK(CLK), .Q(n8825), .QN(n12518)
         );
  DFF_X1 \REGISTERS_reg[9][62]  ( .D(n6474), .CK(CLK), .Q(n8826), .QN(n12519)
         );
  DFF_X1 \REGISTERS_reg[9][61]  ( .D(n6473), .CK(CLK), .Q(n8827), .QN(n12520)
         );
  DFF_X1 \REGISTERS_reg[9][60]  ( .D(n6472), .CK(CLK), .Q(n8828), .QN(n12521)
         );
  DFF_X1 \REGISTERS_reg[11][63]  ( .D(n6347), .CK(CLK), .Q(n8761), .QN(n12646)
         );
  DFF_X1 \REGISTERS_reg[11][62]  ( .D(n6346), .CK(CLK), .Q(n8762), .QN(n12647)
         );
  DFF_X1 \REGISTERS_reg[11][61]  ( .D(n6345), .CK(CLK), .Q(n8763), .QN(n12648)
         );
  DFF_X1 \REGISTERS_reg[11][60]  ( .D(n6344), .CK(CLK), .Q(n8764), .QN(n12649)
         );
  DFF_X1 \REGISTERS_reg[27][63]  ( .D(n5323), .CK(CLK), .Q(n8249), .QN(n13315)
         );
  DFF_X1 \REGISTERS_reg[27][62]  ( .D(n5322), .CK(CLK), .Q(n8250), .QN(n13316)
         );
  DFF_X1 \REGISTERS_reg[27][61]  ( .D(n5321), .CK(CLK), .Q(n8251), .QN(n13317)
         );
  DFF_X1 \REGISTERS_reg[27][60]  ( .D(n5320), .CK(CLK), .Q(n8252), .QN(n13318)
         );
  DFF_X1 \REGISTERS_reg[26][63]  ( .D(n5387), .CK(CLK), .Q(n8569), .QN(n13251)
         );
  DFF_X1 \REGISTERS_reg[26][62]  ( .D(n5386), .CK(CLK), .Q(n8570), .QN(n13252)
         );
  DFF_X1 \REGISTERS_reg[26][61]  ( .D(n5385), .CK(CLK), .Q(n8571), .QN(n13253)
         );
  DFF_X1 \REGISTERS_reg[26][60]  ( .D(n5384), .CK(CLK), .Q(n8572), .QN(n13254)
         );
  DFF_X1 \REGISTERS_reg[8][63]  ( .D(n6539), .CK(CLK), .Q(n8057), .QN(n12454)
         );
  DFF_X1 \REGISTERS_reg[8][62]  ( .D(n6538), .CK(CLK), .Q(n8058), .QN(n12455)
         );
  DFF_X1 \REGISTERS_reg[8][61]  ( .D(n6537), .CK(CLK), .Q(n8059), .QN(n12456)
         );
  DFF_X1 \REGISTERS_reg[8][60]  ( .D(n6536), .CK(CLK), .Q(n8060), .QN(n12457)
         );
  DFF_X1 \REGISTERS_reg[9][59]  ( .D(n6471), .CK(CLK), .Q(n8829), .QN(n12522)
         );
  DFF_X1 \REGISTERS_reg[9][58]  ( .D(n6470), .CK(CLK), .Q(n8830), .QN(n12523)
         );
  DFF_X1 \REGISTERS_reg[9][57]  ( .D(n6469), .CK(CLK), .Q(n8831), .QN(n12524)
         );
  DFF_X1 \REGISTERS_reg[9][56]  ( .D(n6468), .CK(CLK), .Q(n8832), .QN(n12525)
         );
  DFF_X1 \REGISTERS_reg[9][55]  ( .D(n6467), .CK(CLK), .Q(n8833), .QN(n12526)
         );
  DFF_X1 \REGISTERS_reg[9][54]  ( .D(n6466), .CK(CLK), .Q(n8834), .QN(n12527)
         );
  DFF_X1 \REGISTERS_reg[9][53]  ( .D(n6465), .CK(CLK), .Q(n8835), .QN(n12528)
         );
  DFF_X1 \REGISTERS_reg[9][52]  ( .D(n6464), .CK(CLK), .Q(n8836), .QN(n12529)
         );
  DFF_X1 \REGISTERS_reg[9][51]  ( .D(n6463), .CK(CLK), .Q(n8837), .QN(n12530)
         );
  DFF_X1 \REGISTERS_reg[9][50]  ( .D(n6462), .CK(CLK), .Q(n8838), .QN(n12531)
         );
  DFF_X1 \REGISTERS_reg[9][49]  ( .D(n6461), .CK(CLK), .Q(n8839), .QN(n12532)
         );
  DFF_X1 \REGISTERS_reg[9][48]  ( .D(n6460), .CK(CLK), .Q(n8840), .QN(n12533)
         );
  DFF_X1 \REGISTERS_reg[9][47]  ( .D(n6459), .CK(CLK), .Q(n8841), .QN(n12534)
         );
  DFF_X1 \REGISTERS_reg[9][46]  ( .D(n6458), .CK(CLK), .Q(n8842), .QN(n12535)
         );
  DFF_X1 \REGISTERS_reg[9][45]  ( .D(n6457), .CK(CLK), .Q(n8843), .QN(n12536)
         );
  DFF_X1 \REGISTERS_reg[9][44]  ( .D(n6456), .CK(CLK), .Q(n8844), .QN(n12537)
         );
  DFF_X1 \REGISTERS_reg[9][43]  ( .D(n6455), .CK(CLK), .Q(n8845), .QN(n12538)
         );
  DFF_X1 \REGISTERS_reg[9][42]  ( .D(n6454), .CK(CLK), .Q(n8846), .QN(n12539)
         );
  DFF_X1 \REGISTERS_reg[9][41]  ( .D(n6453), .CK(CLK), .Q(n8847), .QN(n12540)
         );
  DFF_X1 \REGISTERS_reg[9][40]  ( .D(n6452), .CK(CLK), .Q(n8848), .QN(n12541)
         );
  DFF_X1 \REGISTERS_reg[9][39]  ( .D(n6451), .CK(CLK), .Q(n8849), .QN(n12542)
         );
  DFF_X1 \REGISTERS_reg[9][38]  ( .D(n6450), .CK(CLK), .Q(n8850), .QN(n12543)
         );
  DFF_X1 \REGISTERS_reg[9][37]  ( .D(n6449), .CK(CLK), .Q(n8851), .QN(n12544)
         );
  DFF_X1 \REGISTERS_reg[9][36]  ( .D(n6448), .CK(CLK), .Q(n8852), .QN(n12545)
         );
  DFF_X1 \REGISTERS_reg[9][35]  ( .D(n6447), .CK(CLK), .Q(n8853), .QN(n12546)
         );
  DFF_X1 \REGISTERS_reg[9][34]  ( .D(n6446), .CK(CLK), .Q(n8854), .QN(n12547)
         );
  DFF_X1 \REGISTERS_reg[9][33]  ( .D(n6445), .CK(CLK), .Q(n8855), .QN(n12548)
         );
  DFF_X1 \REGISTERS_reg[9][32]  ( .D(n6444), .CK(CLK), .Q(n8856), .QN(n12549)
         );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n6443), .CK(CLK), .Q(n8857), .QN(n12550)
         );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n6442), .CK(CLK), .Q(n8858), .QN(n12551)
         );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n6441), .CK(CLK), .Q(n8859), .QN(n12552)
         );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n6440), .CK(CLK), .Q(n8860), .QN(n12553)
         );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n6439), .CK(CLK), .Q(n8861), .QN(n12554)
         );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n6438), .CK(CLK), .Q(n8862), .QN(n12555)
         );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n6437), .CK(CLK), .Q(n8863), .QN(n12556)
         );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n6436), .CK(CLK), .Q(n8864), .QN(n12557)
         );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n6435), .CK(CLK), .Q(n8865), .QN(n12558)
         );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n6434), .CK(CLK), .Q(n8866), .QN(n12559)
         );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n6433), .CK(CLK), .Q(n8867), .QN(n12560)
         );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n6432), .CK(CLK), .Q(n8868), .QN(n12561)
         );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n6431), .CK(CLK), .Q(n8869), .QN(n12562)
         );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n6430), .CK(CLK), .Q(n8870), .QN(n12563)
         );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n6429), .CK(CLK), .Q(n8871), .QN(n12564)
         );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n6428), .CK(CLK), .Q(n8872), .QN(n12565)
         );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n6427), .CK(CLK), .Q(n8873), .QN(n12566)
         );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n6426), .CK(CLK), .Q(n8874), .QN(n12567)
         );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n6425), .CK(CLK), .Q(n8875), .QN(n12568)
         );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n6424), .CK(CLK), .Q(n8876), .QN(n12569)
         );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n6423), .CK(CLK), .Q(n8877), .QN(n12570)
         );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n6422), .CK(CLK), .Q(n8878), .QN(n12571)
         );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n6421), .CK(CLK), .Q(n8879), .QN(n12572)
         );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n6420), .CK(CLK), .Q(n8880), .QN(n12573)
         );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n6419), .CK(CLK), .Q(n8881), .QN(n12574)
         );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n6418), .CK(CLK), .Q(n8882), .QN(n12575)
         );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n6417), .CK(CLK), .Q(n8883), .QN(n12576)
         );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n6416), .CK(CLK), .Q(n8884), .QN(n12577)
         );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n6415), .CK(CLK), .Q(n8885), .QN(n12578)
         );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n6414), .CK(CLK), .Q(n8886), .QN(n12579)
         );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n6413), .CK(CLK), .Q(n8887), .QN(n12580)
         );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n6412), .CK(CLK), .Q(n8888), .QN(n12581)
         );
  DFF_X1 \REGISTERS_reg[11][59]  ( .D(n6343), .CK(CLK), .Q(n8765), .QN(n12650)
         );
  DFF_X1 \REGISTERS_reg[11][58]  ( .D(n6342), .CK(CLK), .Q(n8766), .QN(n12651)
         );
  DFF_X1 \REGISTERS_reg[11][57]  ( .D(n6341), .CK(CLK), .Q(n8767), .QN(n12652)
         );
  DFF_X1 \REGISTERS_reg[11][56]  ( .D(n6340), .CK(CLK), .Q(n8768), .QN(n12653)
         );
  DFF_X1 \REGISTERS_reg[11][55]  ( .D(n6339), .CK(CLK), .Q(n8769), .QN(n12654)
         );
  DFF_X1 \REGISTERS_reg[11][54]  ( .D(n6338), .CK(CLK), .Q(n8770), .QN(n12655)
         );
  DFF_X1 \REGISTERS_reg[11][53]  ( .D(n6337), .CK(CLK), .Q(n8771), .QN(n12656)
         );
  DFF_X1 \REGISTERS_reg[11][52]  ( .D(n6336), .CK(CLK), .Q(n8772), .QN(n12657)
         );
  DFF_X1 \REGISTERS_reg[11][51]  ( .D(n6335), .CK(CLK), .Q(n8773), .QN(n12658)
         );
  DFF_X1 \REGISTERS_reg[11][50]  ( .D(n6334), .CK(CLK), .Q(n8774), .QN(n12659)
         );
  DFF_X1 \REGISTERS_reg[11][49]  ( .D(n6333), .CK(CLK), .Q(n8775), .QN(n12660)
         );
  DFF_X1 \REGISTERS_reg[11][48]  ( .D(n6332), .CK(CLK), .Q(n8776), .QN(n12661)
         );
  DFF_X1 \REGISTERS_reg[11][47]  ( .D(n6331), .CK(CLK), .Q(n8777), .QN(n12662)
         );
  DFF_X1 \REGISTERS_reg[11][46]  ( .D(n6330), .CK(CLK), .Q(n8778), .QN(n12663)
         );
  DFF_X1 \REGISTERS_reg[11][45]  ( .D(n6329), .CK(CLK), .Q(n8779), .QN(n12664)
         );
  DFF_X1 \REGISTERS_reg[11][44]  ( .D(n6328), .CK(CLK), .Q(n8780), .QN(n12665)
         );
  DFF_X1 \REGISTERS_reg[11][43]  ( .D(n6327), .CK(CLK), .Q(n8781), .QN(n12666)
         );
  DFF_X1 \REGISTERS_reg[11][42]  ( .D(n6326), .CK(CLK), .Q(n8782), .QN(n12667)
         );
  DFF_X1 \REGISTERS_reg[11][41]  ( .D(n6325), .CK(CLK), .Q(n8783), .QN(n12668)
         );
  DFF_X1 \REGISTERS_reg[11][40]  ( .D(n6324), .CK(CLK), .Q(n8784), .QN(n12669)
         );
  DFF_X1 \REGISTERS_reg[11][39]  ( .D(n6323), .CK(CLK), .Q(n8785), .QN(n12670)
         );
  DFF_X1 \REGISTERS_reg[11][38]  ( .D(n6322), .CK(CLK), .Q(n8786), .QN(n12671)
         );
  DFF_X1 \REGISTERS_reg[11][37]  ( .D(n6321), .CK(CLK), .Q(n8787), .QN(n12672)
         );
  DFF_X1 \REGISTERS_reg[11][36]  ( .D(n6320), .CK(CLK), .Q(n8788), .QN(n12673)
         );
  DFF_X1 \REGISTERS_reg[11][35]  ( .D(n6319), .CK(CLK), .Q(n8789), .QN(n12674)
         );
  DFF_X1 \REGISTERS_reg[11][34]  ( .D(n6318), .CK(CLK), .Q(n8790), .QN(n12675)
         );
  DFF_X1 \REGISTERS_reg[11][33]  ( .D(n6317), .CK(CLK), .Q(n8791), .QN(n12676)
         );
  DFF_X1 \REGISTERS_reg[11][32]  ( .D(n6316), .CK(CLK), .Q(n8792), .QN(n12677)
         );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n6315), .CK(CLK), .Q(n8793), .QN(n12678)
         );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n6314), .CK(CLK), .Q(n8794), .QN(n12679)
         );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n6313), .CK(CLK), .Q(n8795), .QN(n12680)
         );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n6312), .CK(CLK), .Q(n8796), .QN(n12681)
         );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n6311), .CK(CLK), .Q(n8797), .QN(n12682)
         );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n6310), .CK(CLK), .Q(n8798), .QN(n12683)
         );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n6309), .CK(CLK), .Q(n8799), .QN(n12684)
         );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n6308), .CK(CLK), .Q(n8800), .QN(n12685)
         );
  DFF_X1 \REGISTERS_reg[27][59]  ( .D(n5319), .CK(CLK), .Q(n8253), .QN(n13319)
         );
  DFF_X1 \REGISTERS_reg[27][58]  ( .D(n5318), .CK(CLK), .Q(n8254), .QN(n13320)
         );
  DFF_X1 \REGISTERS_reg[27][57]  ( .D(n5317), .CK(CLK), .Q(n8255), .QN(n13321)
         );
  DFF_X1 \REGISTERS_reg[27][56]  ( .D(n5316), .CK(CLK), .Q(n8256), .QN(n13322)
         );
  DFF_X1 \REGISTERS_reg[27][55]  ( .D(n5315), .CK(CLK), .Q(n8257), .QN(n13323)
         );
  DFF_X1 \REGISTERS_reg[27][54]  ( .D(n5314), .CK(CLK), .Q(n8258), .QN(n13324)
         );
  DFF_X1 \REGISTERS_reg[27][53]  ( .D(n5313), .CK(CLK), .Q(n8259), .QN(n13325)
         );
  DFF_X1 \REGISTERS_reg[27][52]  ( .D(n5312), .CK(CLK), .Q(n8260), .QN(n13326)
         );
  DFF_X1 \REGISTERS_reg[27][51]  ( .D(n5311), .CK(CLK), .Q(n8261), .QN(n13327)
         );
  DFF_X1 \REGISTERS_reg[27][50]  ( .D(n5310), .CK(CLK), .Q(n8262), .QN(n13328)
         );
  DFF_X1 \REGISTERS_reg[27][49]  ( .D(n5309), .CK(CLK), .Q(n8263), .QN(n13329)
         );
  DFF_X1 \REGISTERS_reg[27][48]  ( .D(n5308), .CK(CLK), .Q(n8264), .QN(n13330)
         );
  DFF_X1 \REGISTERS_reg[27][47]  ( .D(n5307), .CK(CLK), .Q(n8265), .QN(n13331)
         );
  DFF_X1 \REGISTERS_reg[27][46]  ( .D(n5306), .CK(CLK), .Q(n8266), .QN(n13332)
         );
  DFF_X1 \REGISTERS_reg[27][45]  ( .D(n5305), .CK(CLK), .Q(n8267), .QN(n13333)
         );
  DFF_X1 \REGISTERS_reg[27][44]  ( .D(n5304), .CK(CLK), .Q(n8268), .QN(n13334)
         );
  DFF_X1 \REGISTERS_reg[27][43]  ( .D(n5303), .CK(CLK), .Q(n8269), .QN(n13335)
         );
  DFF_X1 \REGISTERS_reg[27][42]  ( .D(n5302), .CK(CLK), .Q(n8270), .QN(n13336)
         );
  DFF_X1 \REGISTERS_reg[27][41]  ( .D(n5301), .CK(CLK), .Q(n8271), .QN(n13337)
         );
  DFF_X1 \REGISTERS_reg[27][40]  ( .D(n5300), .CK(CLK), .Q(n8272), .QN(n13338)
         );
  DFF_X1 \REGISTERS_reg[27][39]  ( .D(n5299), .CK(CLK), .Q(n8273), .QN(n13339)
         );
  DFF_X1 \REGISTERS_reg[27][38]  ( .D(n5298), .CK(CLK), .Q(n8274), .QN(n13340)
         );
  DFF_X1 \REGISTERS_reg[27][37]  ( .D(n5297), .CK(CLK), .Q(n8275), .QN(n13341)
         );
  DFF_X1 \REGISTERS_reg[27][36]  ( .D(n5296), .CK(CLK), .Q(n8276), .QN(n13342)
         );
  DFF_X1 \REGISTERS_reg[27][35]  ( .D(n5295), .CK(CLK), .Q(n8277), .QN(n13343)
         );
  DFF_X1 \REGISTERS_reg[27][34]  ( .D(n5294), .CK(CLK), .Q(n8278), .QN(n13344)
         );
  DFF_X1 \REGISTERS_reg[27][33]  ( .D(n5293), .CK(CLK), .Q(n8279), .QN(n13345)
         );
  DFF_X1 \REGISTERS_reg[27][32]  ( .D(n5292), .CK(CLK), .Q(n8280), .QN(n13346)
         );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n5291), .CK(CLK), .Q(n8281), .QN(n13347)
         );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n5290), .CK(CLK), .Q(n8282), .QN(n13348)
         );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n5289), .CK(CLK), .Q(n8283), .QN(n13349)
         );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n5288), .CK(CLK), .Q(n8284), .QN(n13350)
         );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n5287), .CK(CLK), .Q(n8285), .QN(n13351)
         );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n5286), .CK(CLK), .Q(n8286), .QN(n13352)
         );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n5285), .CK(CLK), .Q(n8287), .QN(n13353)
         );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n5284), .CK(CLK), .Q(n8288), .QN(n13354)
         );
  DFF_X1 \REGISTERS_reg[26][59]  ( .D(n5383), .CK(CLK), .Q(n8573), .QN(n13255)
         );
  DFF_X1 \REGISTERS_reg[26][58]  ( .D(n5382), .CK(CLK), .Q(n8574), .QN(n13256)
         );
  DFF_X1 \REGISTERS_reg[26][57]  ( .D(n5381), .CK(CLK), .Q(n8575), .QN(n13257)
         );
  DFF_X1 \REGISTERS_reg[26][56]  ( .D(n5380), .CK(CLK), .Q(n8576), .QN(n13258)
         );
  DFF_X1 \REGISTERS_reg[26][55]  ( .D(n5379), .CK(CLK), .Q(n8577), .QN(n13259)
         );
  DFF_X1 \REGISTERS_reg[26][54]  ( .D(n5378), .CK(CLK), .Q(n8578), .QN(n13260)
         );
  DFF_X1 \REGISTERS_reg[26][53]  ( .D(n5377), .CK(CLK), .Q(n8579), .QN(n13261)
         );
  DFF_X1 \REGISTERS_reg[26][52]  ( .D(n5376), .CK(CLK), .Q(n8580), .QN(n13262)
         );
  DFF_X1 \REGISTERS_reg[26][51]  ( .D(n5375), .CK(CLK), .Q(n8581), .QN(n13263)
         );
  DFF_X1 \REGISTERS_reg[26][50]  ( .D(n5374), .CK(CLK), .Q(n8582), .QN(n13264)
         );
  DFF_X1 \REGISTERS_reg[26][49]  ( .D(n5373), .CK(CLK), .Q(n8583), .QN(n13265)
         );
  DFF_X1 \REGISTERS_reg[26][48]  ( .D(n5372), .CK(CLK), .Q(n8584), .QN(n13266)
         );
  DFF_X1 \REGISTERS_reg[26][47]  ( .D(n5371), .CK(CLK), .Q(n8585), .QN(n13267)
         );
  DFF_X1 \REGISTERS_reg[26][46]  ( .D(n5370), .CK(CLK), .Q(n8586), .QN(n13268)
         );
  DFF_X1 \REGISTERS_reg[26][45]  ( .D(n5369), .CK(CLK), .Q(n8587), .QN(n13269)
         );
  DFF_X1 \REGISTERS_reg[26][44]  ( .D(n5368), .CK(CLK), .Q(n8588), .QN(n13270)
         );
  DFF_X1 \REGISTERS_reg[26][43]  ( .D(n5367), .CK(CLK), .Q(n8589), .QN(n13271)
         );
  DFF_X1 \REGISTERS_reg[26][42]  ( .D(n5366), .CK(CLK), .Q(n8590), .QN(n13272)
         );
  DFF_X1 \REGISTERS_reg[26][41]  ( .D(n5365), .CK(CLK), .Q(n8591), .QN(n13273)
         );
  DFF_X1 \REGISTERS_reg[26][40]  ( .D(n5364), .CK(CLK), .Q(n8592), .QN(n13274)
         );
  DFF_X1 \REGISTERS_reg[26][39]  ( .D(n5363), .CK(CLK), .Q(n8593), .QN(n13275)
         );
  DFF_X1 \REGISTERS_reg[26][38]  ( .D(n5362), .CK(CLK), .Q(n8594), .QN(n13276)
         );
  DFF_X1 \REGISTERS_reg[26][37]  ( .D(n5361), .CK(CLK), .Q(n8595), .QN(n13277)
         );
  DFF_X1 \REGISTERS_reg[26][36]  ( .D(n5360), .CK(CLK), .Q(n8596), .QN(n13278)
         );
  DFF_X1 \REGISTERS_reg[26][35]  ( .D(n5359), .CK(CLK), .Q(n8597), .QN(n13279)
         );
  DFF_X1 \REGISTERS_reg[26][34]  ( .D(n5358), .CK(CLK), .Q(n8598), .QN(n13280)
         );
  DFF_X1 \REGISTERS_reg[26][33]  ( .D(n5357), .CK(CLK), .Q(n8599), .QN(n13281)
         );
  DFF_X1 \REGISTERS_reg[26][32]  ( .D(n5356), .CK(CLK), .Q(n8600), .QN(n13282)
         );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n5355), .CK(CLK), .Q(n8601), .QN(n13283)
         );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n5354), .CK(CLK), .Q(n8602), .QN(n13284)
         );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n5353), .CK(CLK), .Q(n8603), .QN(n13285)
         );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n5352), .CK(CLK), .Q(n8604), .QN(n13286)
         );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n5351), .CK(CLK), .Q(n8605), .QN(n13287)
         );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n5350), .CK(CLK), .Q(n8606), .QN(n13288)
         );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n5349), .CK(CLK), .Q(n8607), .QN(n13289)
         );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n5348), .CK(CLK), .Q(n8608), .QN(n13290)
         );
  DFF_X1 \REGISTERS_reg[8][59]  ( .D(n6535), .CK(CLK), .Q(n8061), .QN(n12458)
         );
  DFF_X1 \REGISTERS_reg[8][58]  ( .D(n6534), .CK(CLK), .Q(n8062), .QN(n12459)
         );
  DFF_X1 \REGISTERS_reg[8][57]  ( .D(n6533), .CK(CLK), .Q(n8063), .QN(n12460)
         );
  DFF_X1 \REGISTERS_reg[8][56]  ( .D(n6532), .CK(CLK), .Q(n8064), .QN(n12461)
         );
  DFF_X1 \REGISTERS_reg[8][55]  ( .D(n6531), .CK(CLK), .Q(n8065), .QN(n12462)
         );
  DFF_X1 \REGISTERS_reg[8][54]  ( .D(n6530), .CK(CLK), .Q(n8066), .QN(n12463)
         );
  DFF_X1 \REGISTERS_reg[8][53]  ( .D(n6529), .CK(CLK), .Q(n8067), .QN(n12464)
         );
  DFF_X1 \REGISTERS_reg[8][52]  ( .D(n6528), .CK(CLK), .Q(n8068), .QN(n12465)
         );
  DFF_X1 \REGISTERS_reg[8][51]  ( .D(n6527), .CK(CLK), .Q(n8069), .QN(n12466)
         );
  DFF_X1 \REGISTERS_reg[8][50]  ( .D(n6526), .CK(CLK), .Q(n8070), .QN(n12467)
         );
  DFF_X1 \REGISTERS_reg[8][49]  ( .D(n6525), .CK(CLK), .Q(n8071), .QN(n12468)
         );
  DFF_X1 \REGISTERS_reg[8][48]  ( .D(n6524), .CK(CLK), .Q(n8072), .QN(n12469)
         );
  DFF_X1 \REGISTERS_reg[8][47]  ( .D(n6523), .CK(CLK), .Q(n8073), .QN(n12470)
         );
  DFF_X1 \REGISTERS_reg[8][46]  ( .D(n6522), .CK(CLK), .Q(n8074), .QN(n12471)
         );
  DFF_X1 \REGISTERS_reg[8][45]  ( .D(n6521), .CK(CLK), .Q(n8075), .QN(n12472)
         );
  DFF_X1 \REGISTERS_reg[8][44]  ( .D(n6520), .CK(CLK), .Q(n8076), .QN(n12473)
         );
  DFF_X1 \REGISTERS_reg[8][43]  ( .D(n6519), .CK(CLK), .Q(n8077), .QN(n12474)
         );
  DFF_X1 \REGISTERS_reg[8][42]  ( .D(n6518), .CK(CLK), .Q(n8078), .QN(n12475)
         );
  DFF_X1 \REGISTERS_reg[8][41]  ( .D(n6517), .CK(CLK), .Q(n8079), .QN(n12476)
         );
  DFF_X1 \REGISTERS_reg[8][40]  ( .D(n6516), .CK(CLK), .Q(n8080), .QN(n12477)
         );
  DFF_X1 \REGISTERS_reg[8][39]  ( .D(n6515), .CK(CLK), .Q(n8081), .QN(n12478)
         );
  DFF_X1 \REGISTERS_reg[8][38]  ( .D(n6514), .CK(CLK), .Q(n8082), .QN(n12479)
         );
  DFF_X1 \REGISTERS_reg[8][37]  ( .D(n6513), .CK(CLK), .Q(n8083), .QN(n12480)
         );
  DFF_X1 \REGISTERS_reg[8][36]  ( .D(n6512), .CK(CLK), .Q(n8084), .QN(n12481)
         );
  DFF_X1 \REGISTERS_reg[8][35]  ( .D(n6511), .CK(CLK), .Q(n8085), .QN(n12482)
         );
  DFF_X1 \REGISTERS_reg[8][34]  ( .D(n6510), .CK(CLK), .Q(n8086), .QN(n12483)
         );
  DFF_X1 \REGISTERS_reg[8][33]  ( .D(n6509), .CK(CLK), .Q(n8087), .QN(n12484)
         );
  DFF_X1 \REGISTERS_reg[8][32]  ( .D(n6508), .CK(CLK), .Q(n8088), .QN(n12485)
         );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n6507), .CK(CLK), .Q(n8089), .QN(n12486)
         );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n6506), .CK(CLK), .Q(n8090), .QN(n12487)
         );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n6505), .CK(CLK), .Q(n8091), .QN(n12488)
         );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n6504), .CK(CLK), .Q(n8092), .QN(n12489)
         );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n6503), .CK(CLK), .Q(n8093), .QN(n12490)
         );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n6502), .CK(CLK), .Q(n8094), .QN(n12491)
         );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n6501), .CK(CLK), .Q(n8095), .QN(n12492)
         );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n6500), .CK(CLK), .Q(n8096), .QN(n12493)
         );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n6307), .CK(CLK), .Q(n8801), .QN(n12686)
         );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n6306), .CK(CLK), .Q(n8802), .QN(n12687)
         );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n6305), .CK(CLK), .Q(n8803), .QN(n12688)
         );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n6304), .CK(CLK), .Q(n8804), .QN(n12689)
         );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n6303), .CK(CLK), .Q(n8805), .QN(n12690)
         );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n6302), .CK(CLK), .Q(n8806), .QN(n12691)
         );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n6301), .CK(CLK), .Q(n8807), .QN(n12692)
         );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n6300), .CK(CLK), .Q(n8808), .QN(n12693)
         );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n6299), .CK(CLK), .Q(n8809), .QN(n12694)
         );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n6298), .CK(CLK), .Q(n8810), .QN(n12695)
         );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n6297), .CK(CLK), .Q(n8811), .QN(n12696)
         );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n6296), .CK(CLK), .Q(n8812), .QN(n12697)
         );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n6295), .CK(CLK), .Q(n8813), .QN(n12698)
         );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n6294), .CK(CLK), .Q(n8814), .QN(n12699)
         );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n6293), .CK(CLK), .Q(n8815), .QN(n12700)
         );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n6292), .CK(CLK), .Q(n8816), .QN(n12701)
         );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n6291), .CK(CLK), .Q(n8817), .QN(n12702)
         );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n6290), .CK(CLK), .Q(n8818), .QN(n12703)
         );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n6289), .CK(CLK), .Q(n8819), .QN(n12704)
         );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n6288), .CK(CLK), .Q(n8820), .QN(n12705)
         );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n6287), .CK(CLK), .Q(n8821), .QN(n12706)
         );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n6286), .CK(CLK), .Q(n8822), .QN(n12707)
         );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n6285), .CK(CLK), .Q(n8823), .QN(n12708)
         );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n6284), .CK(CLK), .Q(n8824), .QN(n12709)
         );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n5283), .CK(CLK), .Q(n8289), .QN(n13355)
         );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n5282), .CK(CLK), .Q(n8290), .QN(n13356)
         );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n5281), .CK(CLK), .Q(n8291), .QN(n13357)
         );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n5280), .CK(CLK), .Q(n8292), .QN(n13358)
         );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n5279), .CK(CLK), .Q(n8293), .QN(n13359)
         );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n5278), .CK(CLK), .Q(n8294), .QN(n13360)
         );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n5277), .CK(CLK), .Q(n8295), .QN(n13361)
         );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n5276), .CK(CLK), .Q(n8296), .QN(n13362)
         );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n5275), .CK(CLK), .Q(n8297), .QN(n13363)
         );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n5274), .CK(CLK), .Q(n8298), .QN(n13364)
         );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n5273), .CK(CLK), .Q(n8299), .QN(n13365)
         );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n5272), .CK(CLK), .Q(n8300), .QN(n13366)
         );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n5271), .CK(CLK), .Q(n8301), .QN(n13367)
         );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n5270), .CK(CLK), .Q(n8302), .QN(n13368)
         );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n5269), .CK(CLK), .Q(n8303), .QN(n13369)
         );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n5268), .CK(CLK), .Q(n8304), .QN(n13370)
         );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n5267), .CK(CLK), .Q(n8305), .QN(n13371)
         );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n5266), .CK(CLK), .Q(n8306), .QN(n13372)
         );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n5265), .CK(CLK), .Q(n8307), .QN(n13373)
         );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n5264), .CK(CLK), .Q(n8308), .QN(n13374)
         );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n5263), .CK(CLK), .Q(n8309), .QN(n13375)
         );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n5262), .CK(CLK), .Q(n8310), .QN(n13376)
         );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n5261), .CK(CLK), .Q(n8311), .QN(n13377)
         );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n5260), .CK(CLK), .Q(n8312), .QN(n13378)
         );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n5347), .CK(CLK), .Q(n8609), .QN(n13291)
         );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n5346), .CK(CLK), .Q(n8610), .QN(n13292)
         );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n5345), .CK(CLK), .Q(n8611), .QN(n13293)
         );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n5344), .CK(CLK), .Q(n8612), .QN(n13294)
         );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n5343), .CK(CLK), .Q(n8613), .QN(n13295)
         );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n5342), .CK(CLK), .Q(n8614), .QN(n13296)
         );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n5341), .CK(CLK), .Q(n8615), .QN(n13297)
         );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n5340), .CK(CLK), .Q(n8616), .QN(n13298)
         );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n5339), .CK(CLK), .Q(n8617), .QN(n13299)
         );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n5338), .CK(CLK), .Q(n8618), .QN(n13300)
         );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n5337), .CK(CLK), .Q(n8619), .QN(n13301)
         );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n5336), .CK(CLK), .Q(n8620), .QN(n13302)
         );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n5335), .CK(CLK), .Q(n8621), .QN(n13303)
         );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n5334), .CK(CLK), .Q(n8622), .QN(n13304)
         );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n5333), .CK(CLK), .Q(n8623), .QN(n13305)
         );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n5332), .CK(CLK), .Q(n8624), .QN(n13306)
         );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n5331), .CK(CLK), .Q(n8625), .QN(n13307)
         );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n5330), .CK(CLK), .Q(n8626), .QN(n13308)
         );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n5329), .CK(CLK), .Q(n8627), .QN(n13309)
         );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n5328), .CK(CLK), .Q(n8628), .QN(n13310)
         );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n5327), .CK(CLK), .Q(n8629), .QN(n13311)
         );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n5326), .CK(CLK), .Q(n8630), .QN(n13312)
         );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n5325), .CK(CLK), .Q(n8631), .QN(n13313)
         );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n5324), .CK(CLK), .Q(n8632), .QN(n13314)
         );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n6499), .CK(CLK), .Q(n8097), .QN(n12494)
         );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n6498), .CK(CLK), .Q(n8098), .QN(n12495)
         );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n6497), .CK(CLK), .Q(n8099), .QN(n12496)
         );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n6496), .CK(CLK), .Q(n8100), .QN(n12497)
         );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n6495), .CK(CLK), .Q(n8101), .QN(n12498)
         );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n6494), .CK(CLK), .Q(n8102), .QN(n12499)
         );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n6493), .CK(CLK), .Q(n8103), .QN(n12500)
         );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n6492), .CK(CLK), .Q(n8104), .QN(n12501)
         );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n6491), .CK(CLK), .Q(n8105), .QN(n12502)
         );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n6490), .CK(CLK), .Q(n8106), .QN(n12503)
         );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n6489), .CK(CLK), .Q(n8107), .QN(n12504)
         );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n6488), .CK(CLK), .Q(n8108), .QN(n12505)
         );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n6487), .CK(CLK), .Q(n8109), .QN(n12506)
         );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n6486), .CK(CLK), .Q(n8110), .QN(n12507)
         );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n6485), .CK(CLK), .Q(n8111), .QN(n12508)
         );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n6484), .CK(CLK), .Q(n8112), .QN(n12509)
         );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n6483), .CK(CLK), .Q(n8113), .QN(n12510)
         );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n6482), .CK(CLK), .Q(n8114), .QN(n12511)
         );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n6481), .CK(CLK), .Q(n8115), .QN(n12512)
         );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n6480), .CK(CLK), .Q(n8116), .QN(n12513)
         );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n6479), .CK(CLK), .Q(n8117), .QN(n12514)
         );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n6478), .CK(CLK), .Q(n8118), .QN(n12515)
         );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n6477), .CK(CLK), .Q(n8119), .QN(n12516)
         );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n6476), .CK(CLK), .Q(n8120), .QN(n12517)
         );
  DFF_X1 \REGISTERS_reg[20][63]  ( .D(n5771), .CK(CLK), .Q(n8185), .QN(n12931)
         );
  DFF_X1 \REGISTERS_reg[20][62]  ( .D(n5770), .CK(CLK), .Q(n8186), .QN(n12932)
         );
  DFF_X1 \REGISTERS_reg[20][61]  ( .D(n5769), .CK(CLK), .Q(n8187), .QN(n12933)
         );
  DFF_X1 \REGISTERS_reg[20][60]  ( .D(n5768), .CK(CLK), .Q(n8188), .QN(n12934)
         );
  DFF_X1 \REGISTERS_reg[17][63]  ( .D(n5963), .CK(CLK), .Q(n8505), .QN(n12867)
         );
  DFF_X1 \REGISTERS_reg[17][62]  ( .D(n5962), .CK(CLK), .Q(n8506), .QN(n12868)
         );
  DFF_X1 \REGISTERS_reg[17][61]  ( .D(n5961), .CK(CLK), .Q(n8507), .QN(n12869)
         );
  DFF_X1 \REGISTERS_reg[17][60]  ( .D(n5960), .CK(CLK), .Q(n8508), .QN(n12870)
         );
  DFF_X1 \REGISTERS_reg[16][63]  ( .D(n6027), .CK(CLK), .Q(n8889), .QN(n12803)
         );
  DFF_X1 \REGISTERS_reg[16][62]  ( .D(n6026), .CK(CLK), .Q(n8890), .QN(n12804)
         );
  DFF_X1 \REGISTERS_reg[16][61]  ( .D(n6025), .CK(CLK), .Q(n8891), .QN(n12805)
         );
  DFF_X1 \REGISTERS_reg[16][60]  ( .D(n6024), .CK(CLK), .Q(n8892), .QN(n12806)
         );
  DFF_X1 \REGISTERS_reg[20][59]  ( .D(n5767), .CK(CLK), .Q(n8189), .QN(n12935)
         );
  DFF_X1 \REGISTERS_reg[20][58]  ( .D(n5766), .CK(CLK), .Q(n8190), .QN(n12936)
         );
  DFF_X1 \REGISTERS_reg[20][57]  ( .D(n5765), .CK(CLK), .Q(n8191), .QN(n12937)
         );
  DFF_X1 \REGISTERS_reg[20][56]  ( .D(n5764), .CK(CLK), .Q(n8192), .QN(n12938)
         );
  DFF_X1 \REGISTERS_reg[20][55]  ( .D(n5763), .CK(CLK), .Q(n8193), .QN(n12939)
         );
  DFF_X1 \REGISTERS_reg[20][54]  ( .D(n5762), .CK(CLK), .Q(n8194), .QN(n12940)
         );
  DFF_X1 \REGISTERS_reg[20][53]  ( .D(n5761), .CK(CLK), .Q(n8195), .QN(n12941)
         );
  DFF_X1 \REGISTERS_reg[20][52]  ( .D(n5760), .CK(CLK), .Q(n8196), .QN(n12942)
         );
  DFF_X1 \REGISTERS_reg[20][51]  ( .D(n5759), .CK(CLK), .Q(n8197), .QN(n12943)
         );
  DFF_X1 \REGISTERS_reg[20][50]  ( .D(n5758), .CK(CLK), .Q(n8198), .QN(n12944)
         );
  DFF_X1 \REGISTERS_reg[20][49]  ( .D(n5757), .CK(CLK), .Q(n8199), .QN(n12945)
         );
  DFF_X1 \REGISTERS_reg[20][48]  ( .D(n5756), .CK(CLK), .Q(n8200), .QN(n12946)
         );
  DFF_X1 \REGISTERS_reg[20][47]  ( .D(n5755), .CK(CLK), .Q(n8201), .QN(n12947)
         );
  DFF_X1 \REGISTERS_reg[20][46]  ( .D(n5754), .CK(CLK), .Q(n8202), .QN(n12948)
         );
  DFF_X1 \REGISTERS_reg[20][45]  ( .D(n5753), .CK(CLK), .Q(n8203), .QN(n12949)
         );
  DFF_X1 \REGISTERS_reg[20][44]  ( .D(n5752), .CK(CLK), .Q(n8204), .QN(n12950)
         );
  DFF_X1 \REGISTERS_reg[20][43]  ( .D(n5751), .CK(CLK), .Q(n8205), .QN(n12951)
         );
  DFF_X1 \REGISTERS_reg[20][42]  ( .D(n5750), .CK(CLK), .Q(n8206), .QN(n12952)
         );
  DFF_X1 \REGISTERS_reg[20][41]  ( .D(n5749), .CK(CLK), .Q(n8207), .QN(n12953)
         );
  DFF_X1 \REGISTERS_reg[20][40]  ( .D(n5748), .CK(CLK), .Q(n8208), .QN(n12954)
         );
  DFF_X1 \REGISTERS_reg[20][39]  ( .D(n5747), .CK(CLK), .Q(n8209), .QN(n12955)
         );
  DFF_X1 \REGISTERS_reg[20][38]  ( .D(n5746), .CK(CLK), .Q(n8210), .QN(n12956)
         );
  DFF_X1 \REGISTERS_reg[20][37]  ( .D(n5745), .CK(CLK), .Q(n8211), .QN(n12957)
         );
  DFF_X1 \REGISTERS_reg[20][36]  ( .D(n5744), .CK(CLK), .Q(n8212), .QN(n12958)
         );
  DFF_X1 \REGISTERS_reg[20][35]  ( .D(n5743), .CK(CLK), .Q(n8213), .QN(n12959)
         );
  DFF_X1 \REGISTERS_reg[20][34]  ( .D(n5742), .CK(CLK), .Q(n8214), .QN(n12960)
         );
  DFF_X1 \REGISTERS_reg[20][33]  ( .D(n5741), .CK(CLK), .Q(n8215), .QN(n12961)
         );
  DFF_X1 \REGISTERS_reg[20][32]  ( .D(n5740), .CK(CLK), .Q(n8216), .QN(n12962)
         );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n5739), .CK(CLK), .Q(n8217), .QN(n12963)
         );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n5738), .CK(CLK), .Q(n8218), .QN(n12964)
         );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n5737), .CK(CLK), .Q(n8219), .QN(n12965)
         );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n5736), .CK(CLK), .Q(n8220), .QN(n12966)
         );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n5735), .CK(CLK), .Q(n8221), .QN(n12967)
         );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n5734), .CK(CLK), .Q(n8222), .QN(n12968)
         );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n5733), .CK(CLK), .Q(n8223), .QN(n12969)
         );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n5732), .CK(CLK), .Q(n8224), .QN(n12970)
         );
  DFF_X1 \REGISTERS_reg[17][59]  ( .D(n5959), .CK(CLK), .Q(n8509), .QN(n12871)
         );
  DFF_X1 \REGISTERS_reg[17][58]  ( .D(n5958), .CK(CLK), .Q(n8510), .QN(n12872)
         );
  DFF_X1 \REGISTERS_reg[17][57]  ( .D(n5957), .CK(CLK), .Q(n8511), .QN(n12873)
         );
  DFF_X1 \REGISTERS_reg[17][56]  ( .D(n5956), .CK(CLK), .Q(n8512), .QN(n12874)
         );
  DFF_X1 \REGISTERS_reg[17][55]  ( .D(n5955), .CK(CLK), .Q(n8513), .QN(n12875)
         );
  DFF_X1 \REGISTERS_reg[17][54]  ( .D(n5954), .CK(CLK), .Q(n8514), .QN(n12876)
         );
  DFF_X1 \REGISTERS_reg[17][53]  ( .D(n5953), .CK(CLK), .Q(n8515), .QN(n12877)
         );
  DFF_X1 \REGISTERS_reg[17][52]  ( .D(n5952), .CK(CLK), .Q(n8516), .QN(n12878)
         );
  DFF_X1 \REGISTERS_reg[17][51]  ( .D(n5951), .CK(CLK), .Q(n8517), .QN(n12879)
         );
  DFF_X1 \REGISTERS_reg[17][50]  ( .D(n5950), .CK(CLK), .Q(n8518), .QN(n12880)
         );
  DFF_X1 \REGISTERS_reg[17][49]  ( .D(n5949), .CK(CLK), .Q(n8519), .QN(n12881)
         );
  DFF_X1 \REGISTERS_reg[17][48]  ( .D(n5948), .CK(CLK), .Q(n8520), .QN(n12882)
         );
  DFF_X1 \REGISTERS_reg[17][47]  ( .D(n5947), .CK(CLK), .Q(n8521), .QN(n12883)
         );
  DFF_X1 \REGISTERS_reg[17][46]  ( .D(n5946), .CK(CLK), .Q(n8522), .QN(n12884)
         );
  DFF_X1 \REGISTERS_reg[17][45]  ( .D(n5945), .CK(CLK), .Q(n8523), .QN(n12885)
         );
  DFF_X1 \REGISTERS_reg[17][44]  ( .D(n5944), .CK(CLK), .Q(n8524), .QN(n12886)
         );
  DFF_X1 \REGISTERS_reg[17][43]  ( .D(n5943), .CK(CLK), .Q(n8525), .QN(n12887)
         );
  DFF_X1 \REGISTERS_reg[17][42]  ( .D(n5942), .CK(CLK), .Q(n8526), .QN(n12888)
         );
  DFF_X1 \REGISTERS_reg[17][41]  ( .D(n5941), .CK(CLK), .Q(n8527), .QN(n12889)
         );
  DFF_X1 \REGISTERS_reg[17][40]  ( .D(n5940), .CK(CLK), .Q(n8528), .QN(n12890)
         );
  DFF_X1 \REGISTERS_reg[17][39]  ( .D(n5939), .CK(CLK), .Q(n8529), .QN(n12891)
         );
  DFF_X1 \REGISTERS_reg[17][38]  ( .D(n5938), .CK(CLK), .Q(n8530), .QN(n12892)
         );
  DFF_X1 \REGISTERS_reg[17][37]  ( .D(n5937), .CK(CLK), .Q(n8531), .QN(n12893)
         );
  DFF_X1 \REGISTERS_reg[17][36]  ( .D(n5936), .CK(CLK), .Q(n8532), .QN(n12894)
         );
  DFF_X1 \REGISTERS_reg[17][35]  ( .D(n5935), .CK(CLK), .Q(n8533), .QN(n12895)
         );
  DFF_X1 \REGISTERS_reg[17][34]  ( .D(n5934), .CK(CLK), .Q(n8534), .QN(n12896)
         );
  DFF_X1 \REGISTERS_reg[17][33]  ( .D(n5933), .CK(CLK), .Q(n8535), .QN(n12897)
         );
  DFF_X1 \REGISTERS_reg[17][32]  ( .D(n5932), .CK(CLK), .Q(n8536), .QN(n12898)
         );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n5931), .CK(CLK), .Q(n8537), .QN(n12899)
         );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n5930), .CK(CLK), .Q(n8538), .QN(n12900)
         );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n5929), .CK(CLK), .Q(n8539), .QN(n12901)
         );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n5928), .CK(CLK), .Q(n8540), .QN(n12902)
         );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n5927), .CK(CLK), .Q(n8541), .QN(n12903)
         );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n5926), .CK(CLK), .Q(n8542), .QN(n12904)
         );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n5925), .CK(CLK), .Q(n8543), .QN(n12905)
         );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n5924), .CK(CLK), .Q(n8544), .QN(n12906)
         );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n5731), .CK(CLK), .Q(n8225), .QN(n12971)
         );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n5730), .CK(CLK), .Q(n8226), .QN(n12972)
         );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n5729), .CK(CLK), .Q(n8227), .QN(n12973)
         );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n5728), .CK(CLK), .Q(n8228), .QN(n12974)
         );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n5727), .CK(CLK), .Q(n8229), .QN(n12975)
         );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n5726), .CK(CLK), .Q(n8230), .QN(n12976)
         );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n5725), .CK(CLK), .Q(n8231), .QN(n12977)
         );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n5724), .CK(CLK), .Q(n8232), .QN(n12978)
         );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n5723), .CK(CLK), .Q(n8233), .QN(n12979)
         );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n5722), .CK(CLK), .Q(n8234), .QN(n12980)
         );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n5721), .CK(CLK), .Q(n8235), .QN(n12981)
         );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n5720), .CK(CLK), .Q(n8236), .QN(n12982)
         );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n5719), .CK(CLK), .Q(n8237), .QN(n12983)
         );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n5718), .CK(CLK), .Q(n8238), .QN(n12984)
         );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n5717), .CK(CLK), .Q(n8239), .QN(n12985)
         );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n5716), .CK(CLK), .Q(n8240), .QN(n12986)
         );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n5715), .CK(CLK), .Q(n8241), .QN(n12987)
         );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n5714), .CK(CLK), .Q(n8242), .QN(n12988)
         );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n5713), .CK(CLK), .Q(n8243), .QN(n12989)
         );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n5712), .CK(CLK), .Q(n8244), .QN(n12990)
         );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n5711), .CK(CLK), .Q(n8245), .QN(n12991)
         );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n5710), .CK(CLK), .Q(n8246), .QN(n12992)
         );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n5709), .CK(CLK), .Q(n8247), .QN(n12993)
         );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n5708), .CK(CLK), .Q(n8248), .QN(n12994)
         );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n5923), .CK(CLK), .Q(n8545), .QN(n12907)
         );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n5922), .CK(CLK), .Q(n8546), .QN(n12908)
         );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n5921), .CK(CLK), .Q(n8547), .QN(n12909)
         );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n5920), .CK(CLK), .Q(n8548), .QN(n12910)
         );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n5919), .CK(CLK), .Q(n8549), .QN(n12911)
         );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n5918), .CK(CLK), .Q(n8550), .QN(n12912)
         );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n5917), .CK(CLK), .Q(n8551), .QN(n12913)
         );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n5916), .CK(CLK), .Q(n8552), .QN(n12914)
         );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n5915), .CK(CLK), .Q(n8553), .QN(n12915)
         );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n5914), .CK(CLK), .Q(n8554), .QN(n12916)
         );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n5913), .CK(CLK), .Q(n8555), .QN(n12917)
         );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n5912), .CK(CLK), .Q(n8556), .QN(n12918)
         );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n5911), .CK(CLK), .Q(n8557), .QN(n12919)
         );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n5910), .CK(CLK), .Q(n8558), .QN(n12920)
         );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n5909), .CK(CLK), .Q(n8559), .QN(n12921)
         );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n5908), .CK(CLK), .Q(n8560), .QN(n12922)
         );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n5907), .CK(CLK), .Q(n8561), .QN(n12923)
         );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n5906), .CK(CLK), .Q(n8562), .QN(n12924)
         );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n5905), .CK(CLK), .Q(n8563), .QN(n12925)
         );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n5904), .CK(CLK), .Q(n8564), .QN(n12926)
         );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n5903), .CK(CLK), .Q(n8565), .QN(n12927)
         );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n5902), .CK(CLK), .Q(n8566), .QN(n12928)
         );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n5901), .CK(CLK), .Q(n8567), .QN(n12929)
         );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n5900), .CK(CLK), .Q(n8568), .QN(n12930)
         );
  DFF_X1 \REGISTERS_reg[16][59]  ( .D(n6023), .CK(CLK), .Q(n8893), .QN(n12807)
         );
  DFF_X1 \REGISTERS_reg[16][58]  ( .D(n6022), .CK(CLK), .Q(n8894), .QN(n12808)
         );
  DFF_X1 \REGISTERS_reg[16][57]  ( .D(n6021), .CK(CLK), .Q(n8895), .QN(n12809)
         );
  DFF_X1 \REGISTERS_reg[16][56]  ( .D(n6020), .CK(CLK), .Q(n8896), .QN(n12810)
         );
  DFF_X1 \REGISTERS_reg[16][55]  ( .D(n6019), .CK(CLK), .Q(n8897), .QN(n12811)
         );
  DFF_X1 \REGISTERS_reg[16][54]  ( .D(n6018), .CK(CLK), .Q(n8898), .QN(n12812)
         );
  DFF_X1 \REGISTERS_reg[16][53]  ( .D(n6017), .CK(CLK), .Q(n8899), .QN(n12813)
         );
  DFF_X1 \REGISTERS_reg[16][52]  ( .D(n6016), .CK(CLK), .Q(n8900), .QN(n12814)
         );
  DFF_X1 \REGISTERS_reg[16][51]  ( .D(n6015), .CK(CLK), .Q(n8901), .QN(n12815)
         );
  DFF_X1 \REGISTERS_reg[16][50]  ( .D(n6014), .CK(CLK), .Q(n8902), .QN(n12816)
         );
  DFF_X1 \REGISTERS_reg[16][49]  ( .D(n6013), .CK(CLK), .Q(n8903), .QN(n12817)
         );
  DFF_X1 \REGISTERS_reg[16][48]  ( .D(n6012), .CK(CLK), .Q(n8904), .QN(n12818)
         );
  DFF_X1 \REGISTERS_reg[16][47]  ( .D(n6011), .CK(CLK), .Q(n8905), .QN(n12819)
         );
  DFF_X1 \REGISTERS_reg[16][46]  ( .D(n6010), .CK(CLK), .Q(n8906), .QN(n12820)
         );
  DFF_X1 \REGISTERS_reg[16][45]  ( .D(n6009), .CK(CLK), .Q(n8907), .QN(n12821)
         );
  DFF_X1 \REGISTERS_reg[16][44]  ( .D(n6008), .CK(CLK), .Q(n8908), .QN(n12822)
         );
  DFF_X1 \REGISTERS_reg[16][43]  ( .D(n6007), .CK(CLK), .Q(n8909), .QN(n12823)
         );
  DFF_X1 \REGISTERS_reg[16][42]  ( .D(n6006), .CK(CLK), .Q(n8910), .QN(n12824)
         );
  DFF_X1 \REGISTERS_reg[16][41]  ( .D(n6005), .CK(CLK), .Q(n8911), .QN(n12825)
         );
  DFF_X1 \REGISTERS_reg[16][40]  ( .D(n6004), .CK(CLK), .Q(n8912), .QN(n12826)
         );
  DFF_X1 \REGISTERS_reg[16][39]  ( .D(n6003), .CK(CLK), .Q(n8913), .QN(n12827)
         );
  DFF_X1 \REGISTERS_reg[16][38]  ( .D(n6002), .CK(CLK), .Q(n8914), .QN(n12828)
         );
  DFF_X1 \REGISTERS_reg[16][37]  ( .D(n6001), .CK(CLK), .Q(n8915), .QN(n12829)
         );
  DFF_X1 \REGISTERS_reg[16][36]  ( .D(n6000), .CK(CLK), .Q(n8916), .QN(n12830)
         );
  DFF_X1 \REGISTERS_reg[16][35]  ( .D(n5999), .CK(CLK), .Q(n8917), .QN(n12831)
         );
  DFF_X1 \REGISTERS_reg[16][34]  ( .D(n5998), .CK(CLK), .Q(n8918), .QN(n12832)
         );
  DFF_X1 \REGISTERS_reg[16][33]  ( .D(n5997), .CK(CLK), .Q(n8919), .QN(n12833)
         );
  DFF_X1 \REGISTERS_reg[16][32]  ( .D(n5996), .CK(CLK), .Q(n8920), .QN(n12834)
         );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n5995), .CK(CLK), .Q(n8921), .QN(n12835)
         );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n5994), .CK(CLK), .Q(n8922), .QN(n12836)
         );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n5993), .CK(CLK), .Q(n8923), .QN(n12837)
         );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n5992), .CK(CLK), .Q(n8924), .QN(n12838)
         );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n5991), .CK(CLK), .Q(n8925), .QN(n12839)
         );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n5990), .CK(CLK), .Q(n8926), .QN(n12840)
         );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n5989), .CK(CLK), .Q(n8927), .QN(n12841)
         );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n5988), .CK(CLK), .Q(n8928), .QN(n12842)
         );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n5987), .CK(CLK), .Q(n8929), .QN(n12843)
         );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n5986), .CK(CLK), .Q(n8930), .QN(n12844)
         );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n5985), .CK(CLK), .Q(n8931), .QN(n12845)
         );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n5984), .CK(CLK), .Q(n8932), .QN(n12846)
         );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n5983), .CK(CLK), .Q(n8933), .QN(n12847)
         );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n5982), .CK(CLK), .Q(n8934), .QN(n12848)
         );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n5981), .CK(CLK), .Q(n8935), .QN(n12849)
         );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n5980), .CK(CLK), .Q(n8936), .QN(n12850)
         );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n5979), .CK(CLK), .Q(n8937), .QN(n12851)
         );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n5978), .CK(CLK), .Q(n8938), .QN(n12852)
         );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n5977), .CK(CLK), .Q(n8939), .QN(n12853)
         );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n5976), .CK(CLK), .Q(n8940), .QN(n12854)
         );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n5975), .CK(CLK), .Q(n8941), .QN(n12855)
         );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n5974), .CK(CLK), .Q(n8942), .QN(n12856)
         );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n5973), .CK(CLK), .Q(n8943), .QN(n12857)
         );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n5972), .CK(CLK), .Q(n8944), .QN(n12858)
         );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n5971), .CK(CLK), .Q(n8945), .QN(n12859)
         );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n5970), .CK(CLK), .Q(n8946), .QN(n12860)
         );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n5969), .CK(CLK), .Q(n8947), .QN(n12861)
         );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n5968), .CK(CLK), .Q(n8948), .QN(n12862)
         );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n5967), .CK(CLK), .Q(n8949), .QN(n12863)
         );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n5966), .CK(CLK), .Q(n8950), .QN(n12864)
         );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n5965), .CK(CLK), .Q(n8951), .QN(n12865)
         );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n5964), .CK(CLK), .Q(n8952), .QN(n12866)
         );
  DFF_X1 \OUT2_reg[63]  ( .D(n4939), .CK(CLK), .Q(OUT2[63]) );
  DFF_X1 \OUT2_reg[62]  ( .D(n4938), .CK(CLK), .Q(OUT2[62]) );
  DFF_X1 \OUT2_reg[61]  ( .D(n4937), .CK(CLK), .Q(OUT2[61]) );
  DFF_X1 \OUT2_reg[60]  ( .D(n4936), .CK(CLK), .Q(OUT2[60]) );
  DFF_X1 \OUT1_reg[63]  ( .D(n5003), .CK(CLK), .Q(OUT1[63]) );
  DFF_X1 \OUT1_reg[62]  ( .D(n5002), .CK(CLK), .Q(OUT1[62]) );
  DFF_X1 \OUT1_reg[61]  ( .D(n5001), .CK(CLK), .Q(OUT1[61]) );
  DFF_X1 \OUT1_reg[60]  ( .D(n5000), .CK(CLK), .Q(OUT1[60]) );
  DFF_X1 \OUT2_reg[59]  ( .D(n4935), .CK(CLK), .Q(OUT2[59]) );
  DFF_X1 \OUT2_reg[58]  ( .D(n4934), .CK(CLK), .Q(OUT2[58]) );
  DFF_X1 \OUT2_reg[57]  ( .D(n4933), .CK(CLK), .Q(OUT2[57]) );
  DFF_X1 \OUT2_reg[56]  ( .D(n4932), .CK(CLK), .Q(OUT2[56]) );
  DFF_X1 \OUT2_reg[55]  ( .D(n4931), .CK(CLK), .Q(OUT2[55]) );
  DFF_X1 \OUT2_reg[54]  ( .D(n4930), .CK(CLK), .Q(OUT2[54]) );
  DFF_X1 \OUT2_reg[53]  ( .D(n4929), .CK(CLK), .Q(OUT2[53]) );
  DFF_X1 \OUT2_reg[52]  ( .D(n4928), .CK(CLK), .Q(OUT2[52]) );
  DFF_X1 \OUT2_reg[51]  ( .D(n4927), .CK(CLK), .Q(OUT2[51]) );
  DFF_X1 \OUT2_reg[50]  ( .D(n4926), .CK(CLK), .Q(OUT2[50]) );
  DFF_X1 \OUT2_reg[49]  ( .D(n4925), .CK(CLK), .Q(OUT2[49]) );
  DFF_X1 \OUT2_reg[48]  ( .D(n4924), .CK(CLK), .Q(OUT2[48]) );
  DFF_X1 \OUT2_reg[47]  ( .D(n4923), .CK(CLK), .Q(OUT2[47]) );
  DFF_X1 \OUT2_reg[46]  ( .D(n4922), .CK(CLK), .Q(OUT2[46]) );
  DFF_X1 \OUT2_reg[45]  ( .D(n4921), .CK(CLK), .Q(OUT2[45]) );
  DFF_X1 \OUT2_reg[44]  ( .D(n4920), .CK(CLK), .Q(OUT2[44]) );
  DFF_X1 \OUT2_reg[43]  ( .D(n4919), .CK(CLK), .Q(OUT2[43]) );
  DFF_X1 \OUT2_reg[42]  ( .D(n4918), .CK(CLK), .Q(OUT2[42]) );
  DFF_X1 \OUT2_reg[41]  ( .D(n4917), .CK(CLK), .Q(OUT2[41]) );
  DFF_X1 \OUT2_reg[40]  ( .D(n4916), .CK(CLK), .Q(OUT2[40]) );
  DFF_X1 \OUT2_reg[39]  ( .D(n4915), .CK(CLK), .Q(OUT2[39]) );
  DFF_X1 \OUT2_reg[38]  ( .D(n4914), .CK(CLK), .Q(OUT2[38]) );
  DFF_X1 \OUT2_reg[37]  ( .D(n4913), .CK(CLK), .Q(OUT2[37]) );
  DFF_X1 \OUT2_reg[36]  ( .D(n4912), .CK(CLK), .Q(OUT2[36]) );
  DFF_X1 \OUT2_reg[35]  ( .D(n4911), .CK(CLK), .Q(OUT2[35]) );
  DFF_X1 \OUT2_reg[34]  ( .D(n4910), .CK(CLK), .Q(OUT2[34]) );
  DFF_X1 \OUT2_reg[33]  ( .D(n4909), .CK(CLK), .Q(OUT2[33]) );
  DFF_X1 \OUT2_reg[32]  ( .D(n4908), .CK(CLK), .Q(OUT2[32]) );
  AND2_X1 U11193 ( .A1(DATAIN[60]), .A2(n17582), .ZN(n16416) );
  AND2_X1 U11194 ( .A1(DATAIN[61]), .A2(n17582), .ZN(n16417) );
  AND2_X1 U11195 ( .A1(DATAIN[62]), .A2(n17582), .ZN(n16418) );
  AND2_X1 U11196 ( .A1(DATAIN[63]), .A2(n17582), .ZN(n16419) );
  AND2_X1 U11197 ( .A1(DATAIN[1]), .A2(n17587), .ZN(n16420) );
  AND2_X1 U11198 ( .A1(DATAIN[2]), .A2(n17587), .ZN(n16421) );
  AND2_X1 U11199 ( .A1(DATAIN[3]), .A2(n17586), .ZN(n16422) );
  AND2_X1 U11200 ( .A1(DATAIN[4]), .A2(n17587), .ZN(n16423) );
  AND2_X1 U11201 ( .A1(DATAIN[5]), .A2(n17586), .ZN(n16424) );
  AND2_X1 U11202 ( .A1(DATAIN[6]), .A2(n17586), .ZN(n16425) );
  AND2_X1 U11203 ( .A1(DATAIN[7]), .A2(n17586), .ZN(n16426) );
  AND2_X1 U11204 ( .A1(DATAIN[8]), .A2(n17586), .ZN(n16427) );
  AND2_X1 U11205 ( .A1(DATAIN[9]), .A2(n17586), .ZN(n16428) );
  AND2_X1 U11206 ( .A1(DATAIN[10]), .A2(n17586), .ZN(n16429) );
  AND2_X1 U11207 ( .A1(DATAIN[11]), .A2(n17586), .ZN(n16430) );
  AND2_X1 U11208 ( .A1(DATAIN[12]), .A2(n17586), .ZN(n16431) );
  AND2_X1 U11209 ( .A1(DATAIN[13]), .A2(n17586), .ZN(n16432) );
  AND2_X1 U11210 ( .A1(DATAIN[14]), .A2(n17586), .ZN(n16433) );
  AND2_X1 U11211 ( .A1(DATAIN[15]), .A2(n17585), .ZN(n16434) );
  AND2_X1 U11212 ( .A1(DATAIN[16]), .A2(n17586), .ZN(n16435) );
  AND2_X1 U11213 ( .A1(DATAIN[17]), .A2(n17585), .ZN(n16436) );
  AND2_X1 U11214 ( .A1(DATAIN[18]), .A2(n17585), .ZN(n16437) );
  AND2_X1 U11215 ( .A1(DATAIN[19]), .A2(n17585), .ZN(n16438) );
  AND2_X1 U11216 ( .A1(DATAIN[20]), .A2(n17585), .ZN(n16439) );
  AND2_X1 U11217 ( .A1(DATAIN[21]), .A2(n17585), .ZN(n16440) );
  AND2_X1 U11218 ( .A1(DATAIN[22]), .A2(n17585), .ZN(n16441) );
  AND2_X1 U11219 ( .A1(DATAIN[23]), .A2(n17584), .ZN(n16442) );
  AND2_X1 U11220 ( .A1(DATAIN[24]), .A2(n17585), .ZN(n16443) );
  AND2_X1 U11221 ( .A1(DATAIN[25]), .A2(n17585), .ZN(n16444) );
  AND2_X1 U11222 ( .A1(DATAIN[26]), .A2(n17585), .ZN(n16445) );
  AND2_X1 U11223 ( .A1(DATAIN[27]), .A2(n17585), .ZN(n16446) );
  AND2_X1 U11224 ( .A1(DATAIN[28]), .A2(n17585), .ZN(n16447) );
  AND2_X1 U11225 ( .A1(DATAIN[29]), .A2(n17584), .ZN(n16448) );
  AND2_X1 U11226 ( .A1(DATAIN[30]), .A2(n17584), .ZN(n16449) );
  AND2_X1 U11227 ( .A1(DATAIN[31]), .A2(n17584), .ZN(n16450) );
  AND2_X1 U11228 ( .A1(DATAIN[32]), .A2(n17584), .ZN(n16451) );
  AND2_X1 U11229 ( .A1(DATAIN[33]), .A2(n17584), .ZN(n16452) );
  AND2_X1 U11230 ( .A1(DATAIN[34]), .A2(n17584), .ZN(n16453) );
  AND2_X1 U11231 ( .A1(DATAIN[35]), .A2(n17584), .ZN(n16454) );
  AND2_X1 U11232 ( .A1(DATAIN[36]), .A2(n17584), .ZN(n16455) );
  AND2_X1 U11233 ( .A1(DATAIN[37]), .A2(n17584), .ZN(n16456) );
  AND2_X1 U11234 ( .A1(DATAIN[38]), .A2(n17584), .ZN(n16457) );
  AND2_X1 U11235 ( .A1(DATAIN[39]), .A2(n17584), .ZN(n16458) );
  AND2_X1 U11236 ( .A1(DATAIN[40]), .A2(n17583), .ZN(n16459) );
  AND2_X1 U11237 ( .A1(DATAIN[41]), .A2(n17583), .ZN(n16460) );
  AND2_X1 U11238 ( .A1(DATAIN[42]), .A2(n17583), .ZN(n16461) );
  AND2_X1 U11239 ( .A1(DATAIN[43]), .A2(n17583), .ZN(n16462) );
  AND2_X1 U11240 ( .A1(DATAIN[44]), .A2(n17583), .ZN(n16463) );
  AND2_X1 U11241 ( .A1(DATAIN[45]), .A2(n17583), .ZN(n16464) );
  AND2_X1 U11242 ( .A1(DATAIN[46]), .A2(n17583), .ZN(n16465) );
  AND2_X1 U11243 ( .A1(DATAIN[47]), .A2(n17583), .ZN(n16466) );
  AND2_X1 U11244 ( .A1(DATAIN[48]), .A2(n17583), .ZN(n16467) );
  AND2_X1 U11245 ( .A1(DATAIN[49]), .A2(n17583), .ZN(n16468) );
  AND2_X1 U11246 ( .A1(DATAIN[50]), .A2(n17583), .ZN(n16469) );
  AND2_X1 U11247 ( .A1(DATAIN[51]), .A2(n17583), .ZN(n16470) );
  AND2_X1 U11248 ( .A1(DATAIN[52]), .A2(n17582), .ZN(n16471) );
  AND2_X1 U11249 ( .A1(DATAIN[53]), .A2(n17582), .ZN(n16472) );
  AND2_X1 U11250 ( .A1(DATAIN[54]), .A2(n17582), .ZN(n16473) );
  AND2_X1 U11251 ( .A1(DATAIN[55]), .A2(n17582), .ZN(n16474) );
  AND2_X1 U11252 ( .A1(DATAIN[56]), .A2(n17582), .ZN(n16475) );
  AND2_X1 U11253 ( .A1(DATAIN[57]), .A2(n17582), .ZN(n16476) );
  AND2_X1 U11254 ( .A1(DATAIN[58]), .A2(n17582), .ZN(n16477) );
  AND2_X1 U11255 ( .A1(DATAIN[59]), .A2(n17582), .ZN(n16478) );
  AND2_X1 U11256 ( .A1(DATAIN[0]), .A2(n17587), .ZN(n16479) );
  INV_X1 U11257 ( .A(n17574), .ZN(n17559) );
  INV_X1 U11258 ( .A(n17574), .ZN(n17560) );
  INV_X1 U11259 ( .A(n17575), .ZN(n17561) );
  INV_X1 U11260 ( .A(n17178), .ZN(n17164) );
  INV_X1 U11261 ( .A(n16939), .ZN(n16925) );
  INV_X1 U11262 ( .A(n16939), .ZN(n16926) );
  INV_X1 U11263 ( .A(n16956), .ZN(n16942) );
  INV_X1 U11264 ( .A(n16956), .ZN(n16943) );
  INV_X1 U11265 ( .A(n17007), .ZN(n16993) );
  INV_X1 U11266 ( .A(n17007), .ZN(n16994) );
  INV_X1 U11267 ( .A(n17024), .ZN(n17010) );
  INV_X1 U11268 ( .A(n17024), .ZN(n17011) );
  INV_X1 U11269 ( .A(n17041), .ZN(n17027) );
  INV_X1 U11270 ( .A(n17041), .ZN(n17028) );
  INV_X1 U11271 ( .A(n17058), .ZN(n17044) );
  INV_X1 U11272 ( .A(n17058), .ZN(n17045) );
  INV_X1 U11273 ( .A(n17109), .ZN(n17095) );
  INV_X1 U11274 ( .A(n17109), .ZN(n17096) );
  INV_X1 U11275 ( .A(n17126), .ZN(n17112) );
  INV_X1 U11276 ( .A(n17126), .ZN(n17113) );
  INV_X1 U11277 ( .A(n17195), .ZN(n17181) );
  INV_X1 U11278 ( .A(n17195), .ZN(n17182) );
  INV_X1 U11279 ( .A(n17212), .ZN(n17198) );
  INV_X1 U11280 ( .A(n17212), .ZN(n17199) );
  INV_X1 U11281 ( .A(n17315), .ZN(n17300) );
  INV_X1 U11282 ( .A(n17315), .ZN(n17301) );
  INV_X1 U11283 ( .A(n17334), .ZN(n17319) );
  INV_X1 U11284 ( .A(n17334), .ZN(n17320) );
  INV_X1 U11285 ( .A(n17353), .ZN(n17338) );
  INV_X1 U11286 ( .A(n17353), .ZN(n17339) );
  INV_X1 U11287 ( .A(n17372), .ZN(n17357) );
  INV_X1 U11288 ( .A(n17372), .ZN(n17358) );
  INV_X1 U11289 ( .A(n17391), .ZN(n17376) );
  INV_X1 U11290 ( .A(n17391), .ZN(n17377) );
  INV_X1 U11291 ( .A(n17410), .ZN(n17395) );
  INV_X1 U11292 ( .A(n17410), .ZN(n17396) );
  INV_X1 U11293 ( .A(n17429), .ZN(n17414) );
  INV_X1 U11294 ( .A(n17429), .ZN(n17415) );
  INV_X1 U11295 ( .A(n17316), .ZN(n17302) );
  INV_X1 U11296 ( .A(n17335), .ZN(n17321) );
  INV_X1 U11297 ( .A(n17354), .ZN(n17340) );
  INV_X1 U11298 ( .A(n17373), .ZN(n17359) );
  INV_X1 U11299 ( .A(n17392), .ZN(n17378) );
  INV_X1 U11300 ( .A(n17411), .ZN(n17397) );
  INV_X1 U11301 ( .A(n17430), .ZN(n17416) );
  INV_X1 U11302 ( .A(n17178), .ZN(n17163) );
  INV_X1 U11303 ( .A(n16905), .ZN(n16891) );
  INV_X1 U11304 ( .A(n16905), .ZN(n16892) );
  INV_X1 U11305 ( .A(n16922), .ZN(n16908) );
  INV_X1 U11306 ( .A(n16922), .ZN(n16909) );
  INV_X1 U11307 ( .A(n16973), .ZN(n16959) );
  INV_X1 U11308 ( .A(n16973), .ZN(n16960) );
  INV_X1 U11309 ( .A(n16990), .ZN(n16976) );
  INV_X1 U11310 ( .A(n16990), .ZN(n16977) );
  INV_X1 U11311 ( .A(n17075), .ZN(n17061) );
  INV_X1 U11312 ( .A(n17075), .ZN(n17062) );
  INV_X1 U11313 ( .A(n17092), .ZN(n17078) );
  INV_X1 U11314 ( .A(n17092), .ZN(n17079) );
  INV_X1 U11315 ( .A(n17143), .ZN(n17129) );
  INV_X1 U11316 ( .A(n17143), .ZN(n17130) );
  INV_X1 U11317 ( .A(n17160), .ZN(n17146) );
  INV_X1 U11318 ( .A(n17160), .ZN(n17147) );
  INV_X1 U11319 ( .A(n17229), .ZN(n17215) );
  INV_X1 U11320 ( .A(n17229), .ZN(n17216) );
  INV_X1 U11321 ( .A(n17246), .ZN(n17232) );
  INV_X1 U11322 ( .A(n17246), .ZN(n17233) );
  INV_X1 U11323 ( .A(n17263), .ZN(n17249) );
  INV_X1 U11324 ( .A(n17263), .ZN(n17250) );
  INV_X1 U11325 ( .A(n17280), .ZN(n17266) );
  INV_X1 U11326 ( .A(n17280), .ZN(n17267) );
  INV_X1 U11327 ( .A(n17297), .ZN(n17283) );
  INV_X1 U11328 ( .A(n17297), .ZN(n17284) );
  BUF_X1 U11329 ( .A(n17576), .Z(n17574) );
  BUF_X1 U11330 ( .A(n17576), .Z(n17562) );
  BUF_X1 U11331 ( .A(n17576), .Z(n17563) );
  BUF_X1 U11332 ( .A(n17576), .Z(n17564) );
  BUF_X1 U11333 ( .A(n17576), .Z(n17565) );
  BUF_X1 U11334 ( .A(n17576), .Z(n17566) );
  BUF_X1 U11335 ( .A(n17576), .Z(n17567) );
  BUF_X1 U11336 ( .A(n17576), .Z(n17568) );
  BUF_X1 U11337 ( .A(n17562), .Z(n17569) );
  BUF_X1 U11338 ( .A(n17563), .Z(n17570) );
  BUF_X1 U11339 ( .A(n17564), .Z(n17571) );
  BUF_X1 U11340 ( .A(n17565), .Z(n17572) );
  BUF_X1 U11341 ( .A(n17566), .Z(n17573) );
  BUF_X1 U11342 ( .A(n17567), .Z(n17575) );
  BUF_X1 U11343 ( .A(n14920), .Z(n16571) );
  BUF_X1 U11344 ( .A(n14920), .Z(n16572) );
  BUF_X1 U11345 ( .A(n14920), .Z(n16573) );
  BUF_X1 U11346 ( .A(n14920), .Z(n16574) );
  BUF_X1 U11347 ( .A(n14920), .Z(n16575) );
  BUF_X1 U11348 ( .A(n13712), .Z(n16776) );
  BUF_X1 U11349 ( .A(n13712), .Z(n16777) );
  BUF_X1 U11350 ( .A(n13712), .Z(n16778) );
  BUF_X1 U11351 ( .A(n13712), .Z(n16779) );
  BUF_X1 U11352 ( .A(n13712), .Z(n16780) );
  BUF_X1 U11353 ( .A(n16906), .Z(n16905) );
  BUF_X1 U11354 ( .A(n16923), .Z(n16922) );
  BUF_X1 U11355 ( .A(n16940), .Z(n16939) );
  BUF_X1 U11356 ( .A(n16957), .Z(n16956) );
  BUF_X1 U11357 ( .A(n16974), .Z(n16973) );
  BUF_X1 U11358 ( .A(n16991), .Z(n16990) );
  BUF_X1 U11359 ( .A(n17008), .Z(n17007) );
  BUF_X1 U11360 ( .A(n17025), .Z(n17024) );
  BUF_X1 U11361 ( .A(n17042), .Z(n17041) );
  BUF_X1 U11362 ( .A(n17059), .Z(n17058) );
  BUF_X1 U11363 ( .A(n17076), .Z(n17075) );
  BUF_X1 U11364 ( .A(n17093), .Z(n17092) );
  BUF_X1 U11365 ( .A(n17110), .Z(n17109) );
  BUF_X1 U11366 ( .A(n17127), .Z(n17126) );
  BUF_X1 U11367 ( .A(n17144), .Z(n17143) );
  BUF_X1 U11368 ( .A(n17161), .Z(n17160) );
  BUF_X1 U11369 ( .A(n17179), .Z(n17177) );
  BUF_X1 U11370 ( .A(n17196), .Z(n17195) );
  BUF_X1 U11371 ( .A(n17213), .Z(n17212) );
  BUF_X1 U11372 ( .A(n17230), .Z(n17229) );
  BUF_X1 U11373 ( .A(n17247), .Z(n17246) );
  BUF_X1 U11374 ( .A(n17264), .Z(n17263) );
  BUF_X1 U11375 ( .A(n17281), .Z(n17280) );
  BUF_X1 U11376 ( .A(n17298), .Z(n17297) );
  BUF_X1 U11377 ( .A(n17317), .Z(n17315) );
  BUF_X1 U11378 ( .A(n17336), .Z(n17334) );
  BUF_X1 U11379 ( .A(n17355), .Z(n17353) );
  BUF_X1 U11380 ( .A(n17374), .Z(n17372) );
  BUF_X1 U11381 ( .A(n17393), .Z(n17391) );
  BUF_X1 U11382 ( .A(n17412), .Z(n17410) );
  BUF_X1 U11383 ( .A(n17431), .Z(n17429) );
  BUF_X1 U11384 ( .A(n16906), .Z(n16893) );
  BUF_X1 U11385 ( .A(n16906), .Z(n16894) );
  BUF_X1 U11386 ( .A(n16906), .Z(n16895) );
  BUF_X1 U11387 ( .A(n16906), .Z(n16896) );
  BUF_X1 U11388 ( .A(n16906), .Z(n16897) );
  BUF_X1 U11389 ( .A(n16906), .Z(n16898) );
  BUF_X1 U11390 ( .A(n16906), .Z(n16899) );
  BUF_X1 U11391 ( .A(n16893), .Z(n16900) );
  BUF_X1 U11392 ( .A(n16894), .Z(n16901) );
  BUF_X1 U11393 ( .A(n16895), .Z(n16902) );
  BUF_X1 U11394 ( .A(n16896), .Z(n16903) );
  BUF_X1 U11395 ( .A(n16897), .Z(n16904) );
  BUF_X1 U11396 ( .A(n16923), .Z(n16910) );
  BUF_X1 U11397 ( .A(n16923), .Z(n16911) );
  BUF_X1 U11398 ( .A(n16923), .Z(n16912) );
  BUF_X1 U11399 ( .A(n16923), .Z(n16913) );
  BUF_X1 U11400 ( .A(n16923), .Z(n16914) );
  BUF_X1 U11401 ( .A(n16923), .Z(n16915) );
  BUF_X1 U11402 ( .A(n16923), .Z(n16916) );
  BUF_X1 U11403 ( .A(n16910), .Z(n16917) );
  BUF_X1 U11404 ( .A(n16911), .Z(n16918) );
  BUF_X1 U11405 ( .A(n16912), .Z(n16919) );
  BUF_X1 U11406 ( .A(n16913), .Z(n16920) );
  BUF_X1 U11407 ( .A(n16914), .Z(n16921) );
  BUF_X1 U11408 ( .A(n16940), .Z(n16927) );
  BUF_X1 U11409 ( .A(n16940), .Z(n16928) );
  BUF_X1 U11410 ( .A(n16940), .Z(n16929) );
  BUF_X1 U11411 ( .A(n16940), .Z(n16930) );
  BUF_X1 U11412 ( .A(n16940), .Z(n16931) );
  BUF_X1 U11413 ( .A(n16940), .Z(n16932) );
  BUF_X1 U11414 ( .A(n16940), .Z(n16933) );
  BUF_X1 U11415 ( .A(n16927), .Z(n16934) );
  BUF_X1 U11416 ( .A(n16928), .Z(n16935) );
  BUF_X1 U11417 ( .A(n16929), .Z(n16936) );
  BUF_X1 U11418 ( .A(n16930), .Z(n16937) );
  BUF_X1 U11419 ( .A(n16931), .Z(n16938) );
  BUF_X1 U11420 ( .A(n16957), .Z(n16944) );
  BUF_X1 U11421 ( .A(n16957), .Z(n16945) );
  BUF_X1 U11422 ( .A(n16957), .Z(n16946) );
  BUF_X1 U11423 ( .A(n16957), .Z(n16947) );
  BUF_X1 U11424 ( .A(n16957), .Z(n16948) );
  BUF_X1 U11425 ( .A(n16957), .Z(n16949) );
  BUF_X1 U11426 ( .A(n16957), .Z(n16950) );
  BUF_X1 U11427 ( .A(n16944), .Z(n16951) );
  BUF_X1 U11428 ( .A(n16945), .Z(n16952) );
  BUF_X1 U11429 ( .A(n16946), .Z(n16953) );
  BUF_X1 U11430 ( .A(n16947), .Z(n16954) );
  BUF_X1 U11431 ( .A(n16948), .Z(n16955) );
  BUF_X1 U11432 ( .A(n16974), .Z(n16961) );
  BUF_X1 U11433 ( .A(n16974), .Z(n16962) );
  BUF_X1 U11434 ( .A(n16974), .Z(n16963) );
  BUF_X1 U11435 ( .A(n16974), .Z(n16964) );
  BUF_X1 U11436 ( .A(n16974), .Z(n16965) );
  BUF_X1 U11437 ( .A(n16974), .Z(n16966) );
  BUF_X1 U11438 ( .A(n16974), .Z(n16967) );
  BUF_X1 U11439 ( .A(n16961), .Z(n16968) );
  BUF_X1 U11440 ( .A(n16962), .Z(n16969) );
  BUF_X1 U11441 ( .A(n16963), .Z(n16970) );
  BUF_X1 U11442 ( .A(n16964), .Z(n16971) );
  BUF_X1 U11443 ( .A(n16965), .Z(n16972) );
  BUF_X1 U11444 ( .A(n16991), .Z(n16978) );
  BUF_X1 U11445 ( .A(n16991), .Z(n16979) );
  BUF_X1 U11446 ( .A(n16991), .Z(n16980) );
  BUF_X1 U11447 ( .A(n16991), .Z(n16981) );
  BUF_X1 U11448 ( .A(n16991), .Z(n16982) );
  BUF_X1 U11449 ( .A(n16991), .Z(n16983) );
  BUF_X1 U11450 ( .A(n16991), .Z(n16984) );
  BUF_X1 U11451 ( .A(n16978), .Z(n16985) );
  BUF_X1 U11452 ( .A(n16979), .Z(n16986) );
  BUF_X1 U11453 ( .A(n16980), .Z(n16987) );
  BUF_X1 U11454 ( .A(n16981), .Z(n16988) );
  BUF_X1 U11455 ( .A(n16982), .Z(n16989) );
  BUF_X1 U11456 ( .A(n17008), .Z(n16995) );
  BUF_X1 U11457 ( .A(n17008), .Z(n16996) );
  BUF_X1 U11458 ( .A(n17008), .Z(n16997) );
  BUF_X1 U11459 ( .A(n17008), .Z(n16998) );
  BUF_X1 U11460 ( .A(n17008), .Z(n16999) );
  BUF_X1 U11461 ( .A(n17008), .Z(n17000) );
  BUF_X1 U11462 ( .A(n17008), .Z(n17001) );
  BUF_X1 U11463 ( .A(n16995), .Z(n17002) );
  BUF_X1 U11464 ( .A(n16996), .Z(n17003) );
  BUF_X1 U11465 ( .A(n16997), .Z(n17004) );
  BUF_X1 U11466 ( .A(n16998), .Z(n17005) );
  BUF_X1 U11467 ( .A(n16999), .Z(n17006) );
  BUF_X1 U11468 ( .A(n17025), .Z(n17012) );
  BUF_X1 U11469 ( .A(n17025), .Z(n17013) );
  BUF_X1 U11470 ( .A(n17025), .Z(n17014) );
  BUF_X1 U11471 ( .A(n17025), .Z(n17015) );
  BUF_X1 U11472 ( .A(n17025), .Z(n17016) );
  BUF_X1 U11473 ( .A(n17025), .Z(n17017) );
  BUF_X1 U11474 ( .A(n17025), .Z(n17018) );
  BUF_X1 U11475 ( .A(n17012), .Z(n17019) );
  BUF_X1 U11476 ( .A(n17013), .Z(n17020) );
  BUF_X1 U11477 ( .A(n17014), .Z(n17021) );
  BUF_X1 U11478 ( .A(n17015), .Z(n17022) );
  BUF_X1 U11479 ( .A(n17016), .Z(n17023) );
  BUF_X1 U11480 ( .A(n17042), .Z(n17029) );
  BUF_X1 U11481 ( .A(n17042), .Z(n17030) );
  BUF_X1 U11482 ( .A(n17042), .Z(n17031) );
  BUF_X1 U11483 ( .A(n17042), .Z(n17032) );
  BUF_X1 U11484 ( .A(n17042), .Z(n17033) );
  BUF_X1 U11485 ( .A(n17042), .Z(n17034) );
  BUF_X1 U11486 ( .A(n17042), .Z(n17035) );
  BUF_X1 U11487 ( .A(n17029), .Z(n17036) );
  BUF_X1 U11488 ( .A(n17030), .Z(n17037) );
  BUF_X1 U11489 ( .A(n17031), .Z(n17038) );
  BUF_X1 U11490 ( .A(n17032), .Z(n17039) );
  BUF_X1 U11491 ( .A(n17033), .Z(n17040) );
  BUF_X1 U11492 ( .A(n17059), .Z(n17046) );
  BUF_X1 U11493 ( .A(n17059), .Z(n17047) );
  BUF_X1 U11494 ( .A(n17059), .Z(n17048) );
  BUF_X1 U11495 ( .A(n17059), .Z(n17049) );
  BUF_X1 U11496 ( .A(n17059), .Z(n17050) );
  BUF_X1 U11497 ( .A(n17059), .Z(n17051) );
  BUF_X1 U11498 ( .A(n17059), .Z(n17052) );
  BUF_X1 U11499 ( .A(n17046), .Z(n17053) );
  BUF_X1 U11500 ( .A(n17047), .Z(n17054) );
  BUF_X1 U11501 ( .A(n17048), .Z(n17055) );
  BUF_X1 U11502 ( .A(n17049), .Z(n17056) );
  BUF_X1 U11503 ( .A(n17050), .Z(n17057) );
  BUF_X1 U11504 ( .A(n17076), .Z(n17063) );
  BUF_X1 U11505 ( .A(n17076), .Z(n17064) );
  BUF_X1 U11506 ( .A(n17076), .Z(n17065) );
  BUF_X1 U11507 ( .A(n17076), .Z(n17066) );
  BUF_X1 U11508 ( .A(n17076), .Z(n17067) );
  BUF_X1 U11509 ( .A(n17076), .Z(n17068) );
  BUF_X1 U11510 ( .A(n17076), .Z(n17069) );
  BUF_X1 U11511 ( .A(n17063), .Z(n17070) );
  BUF_X1 U11512 ( .A(n17064), .Z(n17071) );
  BUF_X1 U11513 ( .A(n17065), .Z(n17072) );
  BUF_X1 U11514 ( .A(n17066), .Z(n17073) );
  BUF_X1 U11515 ( .A(n17067), .Z(n17074) );
  BUF_X1 U11516 ( .A(n17093), .Z(n17080) );
  BUF_X1 U11517 ( .A(n17093), .Z(n17081) );
  BUF_X1 U11518 ( .A(n17093), .Z(n17082) );
  BUF_X1 U11519 ( .A(n17093), .Z(n17083) );
  BUF_X1 U11520 ( .A(n17093), .Z(n17084) );
  BUF_X1 U11521 ( .A(n17093), .Z(n17085) );
  BUF_X1 U11522 ( .A(n17093), .Z(n17086) );
  BUF_X1 U11523 ( .A(n17080), .Z(n17087) );
  BUF_X1 U11524 ( .A(n17081), .Z(n17088) );
  BUF_X1 U11525 ( .A(n17082), .Z(n17089) );
  BUF_X1 U11526 ( .A(n17083), .Z(n17090) );
  BUF_X1 U11527 ( .A(n17084), .Z(n17091) );
  BUF_X1 U11528 ( .A(n17110), .Z(n17097) );
  BUF_X1 U11529 ( .A(n17110), .Z(n17098) );
  BUF_X1 U11530 ( .A(n17110), .Z(n17099) );
  BUF_X1 U11531 ( .A(n17110), .Z(n17100) );
  BUF_X1 U11532 ( .A(n17110), .Z(n17101) );
  BUF_X1 U11533 ( .A(n17110), .Z(n17102) );
  BUF_X1 U11534 ( .A(n17110), .Z(n17103) );
  BUF_X1 U11535 ( .A(n17097), .Z(n17104) );
  BUF_X1 U11536 ( .A(n17098), .Z(n17105) );
  BUF_X1 U11537 ( .A(n17099), .Z(n17106) );
  BUF_X1 U11538 ( .A(n17100), .Z(n17107) );
  BUF_X1 U11539 ( .A(n17101), .Z(n17108) );
  BUF_X1 U11540 ( .A(n17127), .Z(n17114) );
  BUF_X1 U11541 ( .A(n17127), .Z(n17115) );
  BUF_X1 U11542 ( .A(n17127), .Z(n17116) );
  BUF_X1 U11543 ( .A(n17127), .Z(n17117) );
  BUF_X1 U11544 ( .A(n17127), .Z(n17118) );
  BUF_X1 U11545 ( .A(n17127), .Z(n17119) );
  BUF_X1 U11546 ( .A(n17127), .Z(n17120) );
  BUF_X1 U11547 ( .A(n17114), .Z(n17121) );
  BUF_X1 U11548 ( .A(n17115), .Z(n17122) );
  BUF_X1 U11549 ( .A(n17116), .Z(n17123) );
  BUF_X1 U11550 ( .A(n17117), .Z(n17124) );
  BUF_X1 U11551 ( .A(n17118), .Z(n17125) );
  BUF_X1 U11552 ( .A(n17144), .Z(n17131) );
  BUF_X1 U11553 ( .A(n17144), .Z(n17132) );
  BUF_X1 U11554 ( .A(n17144), .Z(n17133) );
  BUF_X1 U11555 ( .A(n17144), .Z(n17134) );
  BUF_X1 U11556 ( .A(n17144), .Z(n17135) );
  BUF_X1 U11557 ( .A(n17144), .Z(n17136) );
  BUF_X1 U11558 ( .A(n17144), .Z(n17137) );
  BUF_X1 U11559 ( .A(n17131), .Z(n17138) );
  BUF_X1 U11560 ( .A(n17132), .Z(n17139) );
  BUF_X1 U11561 ( .A(n17133), .Z(n17140) );
  BUF_X1 U11562 ( .A(n17134), .Z(n17141) );
  BUF_X1 U11563 ( .A(n17135), .Z(n17142) );
  BUF_X1 U11564 ( .A(n17161), .Z(n17148) );
  BUF_X1 U11565 ( .A(n17161), .Z(n17149) );
  BUF_X1 U11566 ( .A(n17161), .Z(n17150) );
  BUF_X1 U11567 ( .A(n17161), .Z(n17151) );
  BUF_X1 U11568 ( .A(n17161), .Z(n17152) );
  BUF_X1 U11569 ( .A(n17161), .Z(n17153) );
  BUF_X1 U11570 ( .A(n17161), .Z(n17154) );
  BUF_X1 U11571 ( .A(n17148), .Z(n17155) );
  BUF_X1 U11572 ( .A(n17149), .Z(n17156) );
  BUF_X1 U11573 ( .A(n17150), .Z(n17157) );
  BUF_X1 U11574 ( .A(n17151), .Z(n17158) );
  BUF_X1 U11575 ( .A(n17152), .Z(n17159) );
  BUF_X1 U11576 ( .A(n17179), .Z(n17165) );
  BUF_X1 U11577 ( .A(n17179), .Z(n17166) );
  BUF_X1 U11578 ( .A(n17179), .Z(n17167) );
  BUF_X1 U11579 ( .A(n17179), .Z(n17168) );
  BUF_X1 U11580 ( .A(n17179), .Z(n17169) );
  BUF_X1 U11581 ( .A(n17179), .Z(n17170) );
  BUF_X1 U11582 ( .A(n17179), .Z(n17171) );
  BUF_X1 U11583 ( .A(n17165), .Z(n17172) );
  BUF_X1 U11584 ( .A(n17166), .Z(n17173) );
  BUF_X1 U11585 ( .A(n17167), .Z(n17174) );
  BUF_X1 U11586 ( .A(n17168), .Z(n17175) );
  BUF_X1 U11587 ( .A(n17169), .Z(n17176) );
  BUF_X1 U11588 ( .A(n17196), .Z(n17183) );
  BUF_X1 U11589 ( .A(n17196), .Z(n17184) );
  BUF_X1 U11590 ( .A(n17196), .Z(n17185) );
  BUF_X1 U11591 ( .A(n17196), .Z(n17186) );
  BUF_X1 U11592 ( .A(n17196), .Z(n17187) );
  BUF_X1 U11593 ( .A(n17196), .Z(n17188) );
  BUF_X1 U11594 ( .A(n17196), .Z(n17189) );
  BUF_X1 U11595 ( .A(n17183), .Z(n17190) );
  BUF_X1 U11596 ( .A(n17184), .Z(n17191) );
  BUF_X1 U11597 ( .A(n17185), .Z(n17192) );
  BUF_X1 U11598 ( .A(n17186), .Z(n17193) );
  BUF_X1 U11599 ( .A(n17187), .Z(n17194) );
  BUF_X1 U11600 ( .A(n17213), .Z(n17200) );
  BUF_X1 U11601 ( .A(n17213), .Z(n17201) );
  BUF_X1 U11602 ( .A(n17213), .Z(n17202) );
  BUF_X1 U11603 ( .A(n17213), .Z(n17203) );
  BUF_X1 U11604 ( .A(n17213), .Z(n17204) );
  BUF_X1 U11605 ( .A(n17213), .Z(n17205) );
  BUF_X1 U11606 ( .A(n17213), .Z(n17206) );
  BUF_X1 U11607 ( .A(n17200), .Z(n17207) );
  BUF_X1 U11608 ( .A(n17201), .Z(n17208) );
  BUF_X1 U11609 ( .A(n17202), .Z(n17209) );
  BUF_X1 U11610 ( .A(n17203), .Z(n17210) );
  BUF_X1 U11611 ( .A(n17204), .Z(n17211) );
  BUF_X1 U11612 ( .A(n17230), .Z(n17217) );
  BUF_X1 U11613 ( .A(n17230), .Z(n17218) );
  BUF_X1 U11614 ( .A(n17230), .Z(n17219) );
  BUF_X1 U11615 ( .A(n17230), .Z(n17220) );
  BUF_X1 U11616 ( .A(n17230), .Z(n17221) );
  BUF_X1 U11617 ( .A(n17230), .Z(n17222) );
  BUF_X1 U11618 ( .A(n17230), .Z(n17223) );
  BUF_X1 U11619 ( .A(n17217), .Z(n17224) );
  BUF_X1 U11620 ( .A(n17218), .Z(n17225) );
  BUF_X1 U11621 ( .A(n17219), .Z(n17226) );
  BUF_X1 U11622 ( .A(n17220), .Z(n17227) );
  BUF_X1 U11623 ( .A(n17221), .Z(n17228) );
  BUF_X1 U11624 ( .A(n17247), .Z(n17234) );
  BUF_X1 U11625 ( .A(n17247), .Z(n17235) );
  BUF_X1 U11626 ( .A(n17247), .Z(n17236) );
  BUF_X1 U11627 ( .A(n17247), .Z(n17237) );
  BUF_X1 U11628 ( .A(n17247), .Z(n17238) );
  BUF_X1 U11629 ( .A(n17247), .Z(n17239) );
  BUF_X1 U11630 ( .A(n17247), .Z(n17240) );
  BUF_X1 U11631 ( .A(n17234), .Z(n17241) );
  BUF_X1 U11632 ( .A(n17235), .Z(n17242) );
  BUF_X1 U11633 ( .A(n17236), .Z(n17243) );
  BUF_X1 U11634 ( .A(n17237), .Z(n17244) );
  BUF_X1 U11635 ( .A(n17238), .Z(n17245) );
  BUF_X1 U11636 ( .A(n17264), .Z(n17251) );
  BUF_X1 U11637 ( .A(n17264), .Z(n17252) );
  BUF_X1 U11638 ( .A(n17264), .Z(n17253) );
  BUF_X1 U11639 ( .A(n17264), .Z(n17254) );
  BUF_X1 U11640 ( .A(n17264), .Z(n17255) );
  BUF_X1 U11641 ( .A(n17264), .Z(n17256) );
  BUF_X1 U11642 ( .A(n17264), .Z(n17257) );
  BUF_X1 U11643 ( .A(n17251), .Z(n17258) );
  BUF_X1 U11644 ( .A(n17252), .Z(n17259) );
  BUF_X1 U11645 ( .A(n17253), .Z(n17260) );
  BUF_X1 U11646 ( .A(n17254), .Z(n17261) );
  BUF_X1 U11647 ( .A(n17255), .Z(n17262) );
  BUF_X1 U11648 ( .A(n17281), .Z(n17268) );
  BUF_X1 U11649 ( .A(n17281), .Z(n17269) );
  BUF_X1 U11650 ( .A(n17281), .Z(n17270) );
  BUF_X1 U11651 ( .A(n17281), .Z(n17271) );
  BUF_X1 U11652 ( .A(n17281), .Z(n17272) );
  BUF_X1 U11653 ( .A(n17281), .Z(n17273) );
  BUF_X1 U11654 ( .A(n17281), .Z(n17274) );
  BUF_X1 U11655 ( .A(n17268), .Z(n17275) );
  BUF_X1 U11656 ( .A(n17269), .Z(n17276) );
  BUF_X1 U11657 ( .A(n17270), .Z(n17277) );
  BUF_X1 U11658 ( .A(n17271), .Z(n17278) );
  BUF_X1 U11659 ( .A(n17272), .Z(n17279) );
  BUF_X1 U11660 ( .A(n17298), .Z(n17285) );
  BUF_X1 U11661 ( .A(n17298), .Z(n17286) );
  BUF_X1 U11662 ( .A(n17298), .Z(n17287) );
  BUF_X1 U11663 ( .A(n17298), .Z(n17288) );
  BUF_X1 U11664 ( .A(n17298), .Z(n17289) );
  BUF_X1 U11665 ( .A(n17298), .Z(n17290) );
  BUF_X1 U11666 ( .A(n17298), .Z(n17291) );
  BUF_X1 U11667 ( .A(n17285), .Z(n17292) );
  BUF_X1 U11668 ( .A(n17286), .Z(n17293) );
  BUF_X1 U11669 ( .A(n17287), .Z(n17294) );
  BUF_X1 U11670 ( .A(n17288), .Z(n17295) );
  BUF_X1 U11671 ( .A(n17289), .Z(n17296) );
  BUF_X1 U11672 ( .A(n17317), .Z(n17303) );
  BUF_X1 U11673 ( .A(n17317), .Z(n17304) );
  BUF_X1 U11674 ( .A(n17317), .Z(n17305) );
  BUF_X1 U11675 ( .A(n17317), .Z(n17306) );
  BUF_X1 U11676 ( .A(n17317), .Z(n17307) );
  BUF_X1 U11677 ( .A(n17317), .Z(n17308) );
  BUF_X1 U11678 ( .A(n17317), .Z(n17309) );
  BUF_X1 U11679 ( .A(n17303), .Z(n17310) );
  BUF_X1 U11680 ( .A(n17304), .Z(n17311) );
  BUF_X1 U11681 ( .A(n17305), .Z(n17312) );
  BUF_X1 U11682 ( .A(n17306), .Z(n17313) );
  BUF_X1 U11683 ( .A(n17307), .Z(n17314) );
  BUF_X1 U11684 ( .A(n17336), .Z(n17322) );
  BUF_X1 U11685 ( .A(n17336), .Z(n17323) );
  BUF_X1 U11686 ( .A(n17336), .Z(n17324) );
  BUF_X1 U11687 ( .A(n17336), .Z(n17325) );
  BUF_X1 U11688 ( .A(n17336), .Z(n17326) );
  BUF_X1 U11689 ( .A(n17336), .Z(n17327) );
  BUF_X1 U11690 ( .A(n17336), .Z(n17328) );
  BUF_X1 U11691 ( .A(n17322), .Z(n17329) );
  BUF_X1 U11692 ( .A(n17323), .Z(n17330) );
  BUF_X1 U11693 ( .A(n17324), .Z(n17331) );
  BUF_X1 U11694 ( .A(n17325), .Z(n17332) );
  BUF_X1 U11695 ( .A(n17326), .Z(n17333) );
  BUF_X1 U11696 ( .A(n17355), .Z(n17341) );
  BUF_X1 U11697 ( .A(n17355), .Z(n17342) );
  BUF_X1 U11698 ( .A(n17355), .Z(n17343) );
  BUF_X1 U11699 ( .A(n17355), .Z(n17344) );
  BUF_X1 U11700 ( .A(n17355), .Z(n17345) );
  BUF_X1 U11701 ( .A(n17355), .Z(n17346) );
  BUF_X1 U11702 ( .A(n17355), .Z(n17347) );
  BUF_X1 U11703 ( .A(n17341), .Z(n17348) );
  BUF_X1 U11704 ( .A(n17342), .Z(n17349) );
  BUF_X1 U11705 ( .A(n17343), .Z(n17350) );
  BUF_X1 U11706 ( .A(n17344), .Z(n17351) );
  BUF_X1 U11707 ( .A(n17345), .Z(n17352) );
  BUF_X1 U11708 ( .A(n17374), .Z(n17360) );
  BUF_X1 U11709 ( .A(n17374), .Z(n17361) );
  BUF_X1 U11710 ( .A(n17374), .Z(n17362) );
  BUF_X1 U11711 ( .A(n17374), .Z(n17363) );
  BUF_X1 U11712 ( .A(n17374), .Z(n17364) );
  BUF_X1 U11713 ( .A(n17374), .Z(n17365) );
  BUF_X1 U11714 ( .A(n17374), .Z(n17366) );
  BUF_X1 U11715 ( .A(n17360), .Z(n17367) );
  BUF_X1 U11716 ( .A(n17361), .Z(n17368) );
  BUF_X1 U11717 ( .A(n17362), .Z(n17369) );
  BUF_X1 U11718 ( .A(n17363), .Z(n17370) );
  BUF_X1 U11719 ( .A(n17364), .Z(n17371) );
  BUF_X1 U11720 ( .A(n17393), .Z(n17379) );
  BUF_X1 U11721 ( .A(n17393), .Z(n17380) );
  BUF_X1 U11722 ( .A(n17393), .Z(n17381) );
  BUF_X1 U11723 ( .A(n17393), .Z(n17382) );
  BUF_X1 U11724 ( .A(n17393), .Z(n17383) );
  BUF_X1 U11725 ( .A(n17393), .Z(n17384) );
  BUF_X1 U11726 ( .A(n17393), .Z(n17385) );
  BUF_X1 U11727 ( .A(n17379), .Z(n17386) );
  BUF_X1 U11728 ( .A(n17380), .Z(n17387) );
  BUF_X1 U11729 ( .A(n17381), .Z(n17388) );
  BUF_X1 U11730 ( .A(n17382), .Z(n17389) );
  BUF_X1 U11731 ( .A(n17383), .Z(n17390) );
  BUF_X1 U11732 ( .A(n17412), .Z(n17398) );
  BUF_X1 U11733 ( .A(n17412), .Z(n17399) );
  BUF_X1 U11734 ( .A(n17412), .Z(n17400) );
  BUF_X1 U11735 ( .A(n17412), .Z(n17401) );
  BUF_X1 U11736 ( .A(n17412), .Z(n17402) );
  BUF_X1 U11737 ( .A(n17412), .Z(n17403) );
  BUF_X1 U11738 ( .A(n17412), .Z(n17404) );
  BUF_X1 U11739 ( .A(n17398), .Z(n17405) );
  BUF_X1 U11740 ( .A(n17399), .Z(n17406) );
  BUF_X1 U11741 ( .A(n17400), .Z(n17407) );
  BUF_X1 U11742 ( .A(n17401), .Z(n17408) );
  BUF_X1 U11743 ( .A(n17402), .Z(n17409) );
  BUF_X1 U11744 ( .A(n17431), .Z(n17417) );
  BUF_X1 U11745 ( .A(n17431), .Z(n17418) );
  BUF_X1 U11746 ( .A(n17431), .Z(n17419) );
  BUF_X1 U11747 ( .A(n17431), .Z(n17420) );
  BUF_X1 U11748 ( .A(n17431), .Z(n17421) );
  BUF_X1 U11749 ( .A(n17431), .Z(n17422) );
  BUF_X1 U11750 ( .A(n17431), .Z(n17423) );
  BUF_X1 U11751 ( .A(n17417), .Z(n17424) );
  BUF_X1 U11752 ( .A(n17418), .Z(n17425) );
  BUF_X1 U11753 ( .A(n17419), .Z(n17426) );
  BUF_X1 U11754 ( .A(n17420), .Z(n17427) );
  BUF_X1 U11755 ( .A(n17421), .Z(n17428) );
  BUF_X1 U11756 ( .A(n17170), .Z(n17178) );
  BUF_X1 U11757 ( .A(n17308), .Z(n17316) );
  BUF_X1 U11758 ( .A(n17327), .Z(n17335) );
  BUF_X1 U11759 ( .A(n17346), .Z(n17354) );
  BUF_X1 U11760 ( .A(n17365), .Z(n17373) );
  BUF_X1 U11761 ( .A(n17384), .Z(n17392) );
  BUF_X1 U11762 ( .A(n17403), .Z(n17411) );
  BUF_X1 U11763 ( .A(n17422), .Z(n17430) );
  INV_X1 U11764 ( .A(n17558), .ZN(n17576) );
  INV_X1 U11765 ( .A(n16479), .ZN(n17432) );
  INV_X1 U11766 ( .A(n16420), .ZN(n17434) );
  INV_X1 U11767 ( .A(n16421), .ZN(n17436) );
  INV_X1 U11768 ( .A(n16422), .ZN(n17438) );
  INV_X1 U11769 ( .A(n16423), .ZN(n17440) );
  INV_X1 U11770 ( .A(n16424), .ZN(n17442) );
  INV_X1 U11771 ( .A(n16425), .ZN(n17444) );
  INV_X1 U11772 ( .A(n16426), .ZN(n17446) );
  INV_X1 U11773 ( .A(n16427), .ZN(n17448) );
  INV_X1 U11774 ( .A(n16428), .ZN(n17450) );
  INV_X1 U11775 ( .A(n16429), .ZN(n17452) );
  INV_X1 U11776 ( .A(n16430), .ZN(n17454) );
  INV_X1 U11777 ( .A(n16431), .ZN(n17456) );
  INV_X1 U11778 ( .A(n16432), .ZN(n17458) );
  INV_X1 U11779 ( .A(n16433), .ZN(n17460) );
  INV_X1 U11780 ( .A(n16434), .ZN(n17462) );
  INV_X1 U11781 ( .A(n16435), .ZN(n17464) );
  INV_X1 U11782 ( .A(n16436), .ZN(n17466) );
  INV_X1 U11783 ( .A(n16437), .ZN(n17468) );
  INV_X1 U11784 ( .A(n16438), .ZN(n17470) );
  INV_X1 U11785 ( .A(n16439), .ZN(n17472) );
  INV_X1 U11786 ( .A(n16440), .ZN(n17474) );
  INV_X1 U11787 ( .A(n16441), .ZN(n17476) );
  INV_X1 U11788 ( .A(n16442), .ZN(n17478) );
  INV_X1 U11789 ( .A(n16443), .ZN(n17480) );
  INV_X1 U11790 ( .A(n16444), .ZN(n17482) );
  INV_X1 U11791 ( .A(n16445), .ZN(n17484) );
  INV_X1 U11792 ( .A(n16446), .ZN(n17486) );
  INV_X1 U11793 ( .A(n16447), .ZN(n17488) );
  INV_X1 U11794 ( .A(n16448), .ZN(n17490) );
  INV_X1 U11795 ( .A(n16449), .ZN(n17492) );
  INV_X1 U11796 ( .A(n16450), .ZN(n17494) );
  INV_X1 U11797 ( .A(n16451), .ZN(n17496) );
  INV_X1 U11798 ( .A(n16452), .ZN(n17498) );
  INV_X1 U11799 ( .A(n16453), .ZN(n17500) );
  INV_X1 U11800 ( .A(n16454), .ZN(n17502) );
  INV_X1 U11801 ( .A(n16455), .ZN(n17504) );
  INV_X1 U11802 ( .A(n16456), .ZN(n17506) );
  INV_X1 U11803 ( .A(n16457), .ZN(n17508) );
  INV_X1 U11804 ( .A(n16458), .ZN(n17510) );
  INV_X1 U11805 ( .A(n16459), .ZN(n17512) );
  INV_X1 U11806 ( .A(n16460), .ZN(n17514) );
  INV_X1 U11807 ( .A(n16461), .ZN(n17516) );
  INV_X1 U11808 ( .A(n16462), .ZN(n17518) );
  INV_X1 U11809 ( .A(n16463), .ZN(n17520) );
  INV_X1 U11810 ( .A(n16464), .ZN(n17522) );
  INV_X1 U11811 ( .A(n16465), .ZN(n17524) );
  INV_X1 U11812 ( .A(n16466), .ZN(n17526) );
  INV_X1 U11813 ( .A(n16467), .ZN(n17528) );
  INV_X1 U11814 ( .A(n16468), .ZN(n17530) );
  INV_X1 U11815 ( .A(n16469), .ZN(n17532) );
  INV_X1 U11816 ( .A(n16470), .ZN(n17534) );
  INV_X1 U11817 ( .A(n16471), .ZN(n17536) );
  INV_X1 U11818 ( .A(n16472), .ZN(n17538) );
  INV_X1 U11819 ( .A(n16473), .ZN(n17540) );
  INV_X1 U11820 ( .A(n16474), .ZN(n17542) );
  INV_X1 U11821 ( .A(n16475), .ZN(n17544) );
  INV_X1 U11822 ( .A(n16476), .ZN(n17546) );
  INV_X1 U11823 ( .A(n16477), .ZN(n17548) );
  INV_X1 U11824 ( .A(n16478), .ZN(n17550) );
  INV_X1 U11825 ( .A(n16416), .ZN(n17552) );
  INV_X1 U11826 ( .A(n16417), .ZN(n17554) );
  INV_X1 U11827 ( .A(n16418), .ZN(n17556) );
  INV_X1 U11828 ( .A(n16419), .ZN(n17577) );
  INV_X1 U11829 ( .A(n16479), .ZN(n17433) );
  INV_X1 U11830 ( .A(n16420), .ZN(n17435) );
  INV_X1 U11831 ( .A(n16421), .ZN(n17437) );
  INV_X1 U11832 ( .A(n16422), .ZN(n17439) );
  INV_X1 U11833 ( .A(n16423), .ZN(n17441) );
  INV_X1 U11834 ( .A(n16424), .ZN(n17443) );
  INV_X1 U11835 ( .A(n16425), .ZN(n17445) );
  INV_X1 U11836 ( .A(n16426), .ZN(n17447) );
  INV_X1 U11837 ( .A(n16427), .ZN(n17449) );
  INV_X1 U11838 ( .A(n16428), .ZN(n17451) );
  INV_X1 U11839 ( .A(n16429), .ZN(n17453) );
  INV_X1 U11840 ( .A(n16430), .ZN(n17455) );
  INV_X1 U11841 ( .A(n16431), .ZN(n17457) );
  INV_X1 U11842 ( .A(n16432), .ZN(n17459) );
  INV_X1 U11843 ( .A(n16433), .ZN(n17461) );
  INV_X1 U11844 ( .A(n16434), .ZN(n17463) );
  INV_X1 U11845 ( .A(n16435), .ZN(n17465) );
  INV_X1 U11846 ( .A(n16436), .ZN(n17467) );
  INV_X1 U11847 ( .A(n16437), .ZN(n17469) );
  INV_X1 U11848 ( .A(n16438), .ZN(n17471) );
  INV_X1 U11849 ( .A(n16439), .ZN(n17473) );
  INV_X1 U11850 ( .A(n16440), .ZN(n17475) );
  INV_X1 U11851 ( .A(n16441), .ZN(n17477) );
  INV_X1 U11852 ( .A(n16442), .ZN(n17479) );
  INV_X1 U11853 ( .A(n16443), .ZN(n17481) );
  INV_X1 U11854 ( .A(n16444), .ZN(n17483) );
  INV_X1 U11855 ( .A(n16445), .ZN(n17485) );
  INV_X1 U11856 ( .A(n16446), .ZN(n17487) );
  INV_X1 U11857 ( .A(n16447), .ZN(n17489) );
  INV_X1 U11858 ( .A(n16448), .ZN(n17491) );
  INV_X1 U11859 ( .A(n16449), .ZN(n17493) );
  INV_X1 U11860 ( .A(n16450), .ZN(n17495) );
  INV_X1 U11861 ( .A(n16451), .ZN(n17497) );
  INV_X1 U11862 ( .A(n16452), .ZN(n17499) );
  INV_X1 U11863 ( .A(n16453), .ZN(n17501) );
  INV_X1 U11864 ( .A(n16454), .ZN(n17503) );
  INV_X1 U11865 ( .A(n16455), .ZN(n17505) );
  INV_X1 U11866 ( .A(n16456), .ZN(n17507) );
  INV_X1 U11867 ( .A(n16457), .ZN(n17509) );
  INV_X1 U11868 ( .A(n16458), .ZN(n17511) );
  INV_X1 U11869 ( .A(n16459), .ZN(n17513) );
  INV_X1 U11870 ( .A(n16460), .ZN(n17515) );
  INV_X1 U11871 ( .A(n16461), .ZN(n17517) );
  INV_X1 U11872 ( .A(n16462), .ZN(n17519) );
  INV_X1 U11873 ( .A(n16463), .ZN(n17521) );
  INV_X1 U11874 ( .A(n16464), .ZN(n17523) );
  INV_X1 U11875 ( .A(n16465), .ZN(n17525) );
  INV_X1 U11876 ( .A(n16466), .ZN(n17527) );
  INV_X1 U11877 ( .A(n16467), .ZN(n17529) );
  INV_X1 U11878 ( .A(n16468), .ZN(n17531) );
  INV_X1 U11879 ( .A(n16469), .ZN(n17533) );
  INV_X1 U11880 ( .A(n16470), .ZN(n17535) );
  INV_X1 U11881 ( .A(n16471), .ZN(n17537) );
  INV_X1 U11882 ( .A(n16472), .ZN(n17539) );
  INV_X1 U11883 ( .A(n16473), .ZN(n17541) );
  INV_X1 U11884 ( .A(n16474), .ZN(n17543) );
  INV_X1 U11885 ( .A(n16475), .ZN(n17545) );
  INV_X1 U11886 ( .A(n16476), .ZN(n17547) );
  INV_X1 U11887 ( .A(n16477), .ZN(n17549) );
  INV_X1 U11888 ( .A(n16478), .ZN(n17551) );
  INV_X1 U11889 ( .A(n16416), .ZN(n17553) );
  INV_X1 U11890 ( .A(n16417), .ZN(n17555) );
  INV_X1 U11891 ( .A(n16418), .ZN(n17557) );
  INV_X1 U11892 ( .A(n16419), .ZN(n17578) );
  BUF_X1 U11893 ( .A(n14910), .Z(n16601) );
  BUF_X1 U11894 ( .A(n14895), .Z(n16673) );
  BUF_X1 U11895 ( .A(n14900), .Z(n16649) );
  BUF_X1 U11896 ( .A(n14905), .Z(n16625) );
  BUF_X1 U11897 ( .A(n14935), .Z(n16500) );
  BUF_X1 U11898 ( .A(n14930), .Z(n16524) );
  BUF_X1 U11899 ( .A(n14910), .Z(n16602) );
  BUF_X1 U11900 ( .A(n14895), .Z(n16674) );
  BUF_X1 U11901 ( .A(n14900), .Z(n16650) );
  BUF_X1 U11902 ( .A(n14905), .Z(n16626) );
  BUF_X1 U11903 ( .A(n14935), .Z(n16501) );
  BUF_X1 U11904 ( .A(n14930), .Z(n16525) );
  BUF_X1 U11905 ( .A(n14910), .Z(n16603) );
  BUF_X1 U11906 ( .A(n14895), .Z(n16675) );
  BUF_X1 U11907 ( .A(n14900), .Z(n16651) );
  BUF_X1 U11908 ( .A(n14905), .Z(n16627) );
  BUF_X1 U11909 ( .A(n14935), .Z(n16502) );
  BUF_X1 U11910 ( .A(n14930), .Z(n16526) );
  BUF_X1 U11911 ( .A(n14910), .Z(n16604) );
  BUF_X1 U11912 ( .A(n14895), .Z(n16676) );
  BUF_X1 U11913 ( .A(n14900), .Z(n16652) );
  BUF_X1 U11914 ( .A(n14905), .Z(n16628) );
  BUF_X1 U11915 ( .A(n14935), .Z(n16503) );
  BUF_X1 U11916 ( .A(n14930), .Z(n16527) );
  BUF_X1 U11917 ( .A(n13702), .Z(n16806) );
  BUF_X1 U11918 ( .A(n13687), .Z(n16878) );
  BUF_X1 U11919 ( .A(n13692), .Z(n16854) );
  BUF_X1 U11920 ( .A(n13697), .Z(n16830) );
  BUF_X1 U11921 ( .A(n13727), .Z(n16705) );
  BUF_X1 U11922 ( .A(n13722), .Z(n16729) );
  BUF_X1 U11923 ( .A(n13702), .Z(n16807) );
  BUF_X1 U11924 ( .A(n13687), .Z(n16879) );
  BUF_X1 U11925 ( .A(n13692), .Z(n16855) );
  BUF_X1 U11926 ( .A(n13697), .Z(n16831) );
  BUF_X1 U11927 ( .A(n13727), .Z(n16706) );
  BUF_X1 U11928 ( .A(n13722), .Z(n16730) );
  BUF_X1 U11929 ( .A(n13702), .Z(n16808) );
  BUF_X1 U11930 ( .A(n13687), .Z(n16880) );
  BUF_X1 U11931 ( .A(n13692), .Z(n16856) );
  BUF_X1 U11932 ( .A(n13697), .Z(n16832) );
  BUF_X1 U11933 ( .A(n13727), .Z(n16707) );
  BUF_X1 U11934 ( .A(n13722), .Z(n16731) );
  BUF_X1 U11935 ( .A(n13702), .Z(n16809) );
  BUF_X1 U11936 ( .A(n13687), .Z(n16881) );
  BUF_X1 U11937 ( .A(n13692), .Z(n16857) );
  BUF_X1 U11938 ( .A(n13697), .Z(n16833) );
  BUF_X1 U11939 ( .A(n13727), .Z(n16708) );
  BUF_X1 U11940 ( .A(n13722), .Z(n16732) );
  BUF_X1 U11941 ( .A(n14909), .Z(n16607) );
  BUF_X1 U11942 ( .A(n14894), .Z(n16679) );
  BUF_X1 U11943 ( .A(n14899), .Z(n16655) );
  BUF_X1 U11944 ( .A(n14904), .Z(n16631) );
  BUF_X1 U11945 ( .A(n14934), .Z(n16506) );
  BUF_X1 U11946 ( .A(n14929), .Z(n16530) );
  BUF_X1 U11947 ( .A(n14909), .Z(n16608) );
  BUF_X1 U11948 ( .A(n14894), .Z(n16680) );
  BUF_X1 U11949 ( .A(n14899), .Z(n16656) );
  BUF_X1 U11950 ( .A(n14904), .Z(n16632) );
  BUF_X1 U11951 ( .A(n14934), .Z(n16507) );
  BUF_X1 U11952 ( .A(n14929), .Z(n16531) );
  BUF_X1 U11953 ( .A(n14909), .Z(n16609) );
  BUF_X1 U11954 ( .A(n14894), .Z(n16681) );
  BUF_X1 U11955 ( .A(n14899), .Z(n16657) );
  BUF_X1 U11956 ( .A(n14904), .Z(n16633) );
  BUF_X1 U11957 ( .A(n14934), .Z(n16508) );
  BUF_X1 U11958 ( .A(n14929), .Z(n16532) );
  BUF_X1 U11959 ( .A(n14909), .Z(n16610) );
  BUF_X1 U11960 ( .A(n14894), .Z(n16682) );
  BUF_X1 U11961 ( .A(n14899), .Z(n16658) );
  BUF_X1 U11962 ( .A(n14904), .Z(n16634) );
  BUF_X1 U11963 ( .A(n14934), .Z(n16509) );
  BUF_X1 U11964 ( .A(n14929), .Z(n16533) );
  BUF_X1 U11965 ( .A(n13701), .Z(n16812) );
  BUF_X1 U11966 ( .A(n13686), .Z(n16884) );
  BUF_X1 U11967 ( .A(n13691), .Z(n16860) );
  BUF_X1 U11968 ( .A(n13696), .Z(n16836) );
  BUF_X1 U11969 ( .A(n13726), .Z(n16711) );
  BUF_X1 U11970 ( .A(n13721), .Z(n16735) );
  BUF_X1 U11971 ( .A(n13701), .Z(n16813) );
  BUF_X1 U11972 ( .A(n13686), .Z(n16885) );
  BUF_X1 U11973 ( .A(n13691), .Z(n16861) );
  BUF_X1 U11974 ( .A(n13696), .Z(n16837) );
  BUF_X1 U11975 ( .A(n13726), .Z(n16712) );
  BUF_X1 U11976 ( .A(n13721), .Z(n16736) );
  BUF_X1 U11977 ( .A(n13701), .Z(n16814) );
  BUF_X1 U11978 ( .A(n13686), .Z(n16886) );
  BUF_X1 U11979 ( .A(n13691), .Z(n16862) );
  BUF_X1 U11980 ( .A(n13696), .Z(n16838) );
  BUF_X1 U11981 ( .A(n13726), .Z(n16713) );
  BUF_X1 U11982 ( .A(n13721), .Z(n16737) );
  BUF_X1 U11983 ( .A(n13701), .Z(n16815) );
  BUF_X1 U11984 ( .A(n13686), .Z(n16887) );
  BUF_X1 U11985 ( .A(n13691), .Z(n16863) );
  BUF_X1 U11986 ( .A(n13696), .Z(n16839) );
  BUF_X1 U11987 ( .A(n13726), .Z(n16714) );
  BUF_X1 U11988 ( .A(n13721), .Z(n16738) );
  BUF_X1 U11989 ( .A(n14912), .Z(n16595) );
  BUF_X1 U11990 ( .A(n14937), .Z(n16494) );
  BUF_X1 U11991 ( .A(n14912), .Z(n16596) );
  BUF_X1 U11992 ( .A(n14937), .Z(n16495) );
  BUF_X1 U11993 ( .A(n14912), .Z(n16597) );
  BUF_X1 U11994 ( .A(n14937), .Z(n16496) );
  BUF_X1 U11995 ( .A(n14912), .Z(n16598) );
  BUF_X1 U11996 ( .A(n14937), .Z(n16497) );
  BUF_X1 U11997 ( .A(n14912), .Z(n16599) );
  BUF_X1 U11998 ( .A(n14937), .Z(n16498) );
  BUF_X1 U11999 ( .A(n13704), .Z(n16800) );
  BUF_X1 U12000 ( .A(n13729), .Z(n16699) );
  BUF_X1 U12001 ( .A(n13704), .Z(n16801) );
  BUF_X1 U12002 ( .A(n13729), .Z(n16700) );
  BUF_X1 U12003 ( .A(n13704), .Z(n16802) );
  BUF_X1 U12004 ( .A(n13729), .Z(n16701) );
  BUF_X1 U12005 ( .A(n13704), .Z(n16803) );
  BUF_X1 U12006 ( .A(n13729), .Z(n16702) );
  BUF_X1 U12007 ( .A(n13704), .Z(n16804) );
  BUF_X1 U12008 ( .A(n13729), .Z(n16703) );
  BUF_X1 U12009 ( .A(n14932), .Z(n16522) );
  BUF_X1 U12010 ( .A(n14932), .Z(n16521) );
  BUF_X1 U12011 ( .A(n14932), .Z(n16520) );
  BUF_X1 U12012 ( .A(n14932), .Z(n16519) );
  BUF_X1 U12013 ( .A(n14897), .Z(n16667) );
  BUF_X1 U12014 ( .A(n14902), .Z(n16643) );
  BUF_X1 U12015 ( .A(n14907), .Z(n16619) );
  BUF_X1 U12016 ( .A(n14897), .Z(n16668) );
  BUF_X1 U12017 ( .A(n14902), .Z(n16644) );
  BUF_X1 U12018 ( .A(n14907), .Z(n16620) );
  BUF_X1 U12019 ( .A(n14897), .Z(n16669) );
  BUF_X1 U12020 ( .A(n14902), .Z(n16645) );
  BUF_X1 U12021 ( .A(n14907), .Z(n16621) );
  BUF_X1 U12022 ( .A(n14897), .Z(n16670) );
  BUF_X1 U12023 ( .A(n14902), .Z(n16646) );
  BUF_X1 U12024 ( .A(n14907), .Z(n16622) );
  BUF_X1 U12025 ( .A(n14897), .Z(n16671) );
  BUF_X1 U12026 ( .A(n14902), .Z(n16647) );
  BUF_X1 U12027 ( .A(n14907), .Z(n16623) );
  BUF_X1 U12028 ( .A(n13689), .Z(n16872) );
  BUF_X1 U12029 ( .A(n13694), .Z(n16848) );
  BUF_X1 U12030 ( .A(n13699), .Z(n16824) );
  BUF_X1 U12031 ( .A(n13689), .Z(n16873) );
  BUF_X1 U12032 ( .A(n13694), .Z(n16849) );
  BUF_X1 U12033 ( .A(n13699), .Z(n16825) );
  BUF_X1 U12034 ( .A(n13689), .Z(n16874) );
  BUF_X1 U12035 ( .A(n13694), .Z(n16850) );
  BUF_X1 U12036 ( .A(n13699), .Z(n16826) );
  BUF_X1 U12037 ( .A(n13689), .Z(n16875) );
  BUF_X1 U12038 ( .A(n13694), .Z(n16851) );
  BUF_X1 U12039 ( .A(n13699), .Z(n16827) );
  BUF_X1 U12040 ( .A(n13689), .Z(n16876) );
  BUF_X1 U12041 ( .A(n13694), .Z(n16852) );
  BUF_X1 U12042 ( .A(n13699), .Z(n16828) );
  BUF_X1 U12043 ( .A(n14922), .Z(n16565) );
  BUF_X1 U12044 ( .A(n14927), .Z(n16546) );
  BUF_X1 U12045 ( .A(n14922), .Z(n16566) );
  BUF_X1 U12046 ( .A(n14927), .Z(n16545) );
  BUF_X1 U12047 ( .A(n14922), .Z(n16567) );
  BUF_X1 U12048 ( .A(n14927), .Z(n16544) );
  BUF_X1 U12049 ( .A(n14922), .Z(n16568) );
  BUF_X1 U12050 ( .A(n14927), .Z(n16543) );
  BUF_X1 U12051 ( .A(n14922), .Z(n16569) );
  BUF_X1 U12052 ( .A(n14927), .Z(n16542) );
  BUF_X1 U12053 ( .A(n13714), .Z(n16770) );
  BUF_X1 U12054 ( .A(n13724), .Z(n16723) );
  BUF_X1 U12055 ( .A(n13719), .Z(n16747) );
  BUF_X1 U12056 ( .A(n13714), .Z(n16771) );
  BUF_X1 U12057 ( .A(n13724), .Z(n16724) );
  BUF_X1 U12058 ( .A(n13719), .Z(n16748) );
  BUF_X1 U12059 ( .A(n13714), .Z(n16772) );
  BUF_X1 U12060 ( .A(n13724), .Z(n16725) );
  BUF_X1 U12061 ( .A(n13719), .Z(n16749) );
  BUF_X1 U12062 ( .A(n13714), .Z(n16773) );
  BUF_X1 U12063 ( .A(n13724), .Z(n16726) );
  BUF_X1 U12064 ( .A(n13719), .Z(n16750) );
  BUF_X1 U12065 ( .A(n13714), .Z(n16774) );
  BUF_X1 U12066 ( .A(n13719), .Z(n16751) );
  BUF_X1 U12067 ( .A(n13724), .Z(n16727) );
  BUF_X1 U12068 ( .A(n14924), .Z(n16555) );
  BUF_X1 U12069 ( .A(n14919), .Z(n16578) );
  BUF_X1 U12070 ( .A(n14924), .Z(n16556) );
  BUF_X1 U12071 ( .A(n14919), .Z(n16579) );
  BUF_X1 U12072 ( .A(n14924), .Z(n16557) );
  BUF_X1 U12073 ( .A(n14919), .Z(n16580) );
  BUF_X1 U12074 ( .A(n14924), .Z(n16558) );
  BUF_X1 U12075 ( .A(n14919), .Z(n16581) );
  BUF_X1 U12076 ( .A(n13711), .Z(n16783) );
  BUF_X1 U12077 ( .A(n13716), .Z(n16760) );
  BUF_X1 U12078 ( .A(n13711), .Z(n16784) );
  BUF_X1 U12079 ( .A(n13716), .Z(n16761) );
  BUF_X1 U12080 ( .A(n13711), .Z(n16785) );
  BUF_X1 U12081 ( .A(n13716), .Z(n16762) );
  BUF_X1 U12082 ( .A(n13711), .Z(n16786) );
  BUF_X1 U12083 ( .A(n13716), .Z(n16763) );
  BUF_X1 U12084 ( .A(n14913), .Z(n16589) );
  BUF_X1 U12085 ( .A(n14938), .Z(n16488) );
  BUF_X1 U12086 ( .A(n14913), .Z(n16590) );
  BUF_X1 U12087 ( .A(n14938), .Z(n16489) );
  BUF_X1 U12088 ( .A(n14913), .Z(n16591) );
  BUF_X1 U12089 ( .A(n14938), .Z(n16490) );
  BUF_X1 U12090 ( .A(n14913), .Z(n16592) );
  BUF_X1 U12091 ( .A(n14938), .Z(n16491) );
  BUF_X1 U12092 ( .A(n14913), .Z(n16593) );
  BUF_X1 U12093 ( .A(n14938), .Z(n16492) );
  BUF_X1 U12094 ( .A(n13705), .Z(n16794) );
  BUF_X1 U12095 ( .A(n13730), .Z(n16693) );
  BUF_X1 U12096 ( .A(n13705), .Z(n16795) );
  BUF_X1 U12097 ( .A(n13730), .Z(n16694) );
  BUF_X1 U12098 ( .A(n13705), .Z(n16796) );
  BUF_X1 U12099 ( .A(n13730), .Z(n16695) );
  BUF_X1 U12100 ( .A(n13705), .Z(n16797) );
  BUF_X1 U12101 ( .A(n13730), .Z(n16696) );
  BUF_X1 U12102 ( .A(n13705), .Z(n16798) );
  BUF_X1 U12103 ( .A(n13730), .Z(n16697) );
  BUF_X1 U12104 ( .A(n14928), .Z(n16536) );
  BUF_X1 U12105 ( .A(n14933), .Z(n16512) );
  BUF_X1 U12106 ( .A(n13720), .Z(n16741) );
  BUF_X1 U12107 ( .A(n13720), .Z(n16742) );
  BUF_X1 U12108 ( .A(n13720), .Z(n16743) );
  BUF_X1 U12109 ( .A(n13720), .Z(n16744) );
  BUF_X1 U12110 ( .A(n13720), .Z(n16745) );
  BUF_X1 U12111 ( .A(n14898), .Z(n16661) );
  BUF_X1 U12112 ( .A(n14903), .Z(n16637) );
  BUF_X1 U12113 ( .A(n14908), .Z(n16613) );
  BUF_X1 U12114 ( .A(n14898), .Z(n16662) );
  BUF_X1 U12115 ( .A(n14903), .Z(n16638) );
  BUF_X1 U12116 ( .A(n14908), .Z(n16614) );
  BUF_X1 U12117 ( .A(n14898), .Z(n16663) );
  BUF_X1 U12118 ( .A(n14903), .Z(n16639) );
  BUF_X1 U12119 ( .A(n14908), .Z(n16615) );
  BUF_X1 U12120 ( .A(n14898), .Z(n16664) );
  BUF_X1 U12121 ( .A(n14903), .Z(n16640) );
  BUF_X1 U12122 ( .A(n14908), .Z(n16616) );
  BUF_X1 U12123 ( .A(n14898), .Z(n16665) );
  BUF_X1 U12124 ( .A(n14903), .Z(n16641) );
  BUF_X1 U12125 ( .A(n14908), .Z(n16617) );
  BUF_X1 U12126 ( .A(n13690), .Z(n16866) );
  BUF_X1 U12127 ( .A(n13695), .Z(n16842) );
  BUF_X1 U12128 ( .A(n13700), .Z(n16818) );
  BUF_X1 U12129 ( .A(n13690), .Z(n16867) );
  BUF_X1 U12130 ( .A(n13695), .Z(n16843) );
  BUF_X1 U12131 ( .A(n13700), .Z(n16819) );
  BUF_X1 U12132 ( .A(n13690), .Z(n16868) );
  BUF_X1 U12133 ( .A(n13695), .Z(n16844) );
  BUF_X1 U12134 ( .A(n13700), .Z(n16820) );
  BUF_X1 U12135 ( .A(n13690), .Z(n16869) );
  BUF_X1 U12136 ( .A(n13695), .Z(n16845) );
  BUF_X1 U12137 ( .A(n13700), .Z(n16821) );
  BUF_X1 U12138 ( .A(n13690), .Z(n16870) );
  BUF_X1 U12139 ( .A(n13695), .Z(n16846) );
  BUF_X1 U12140 ( .A(n13700), .Z(n16822) );
  BUF_X1 U12141 ( .A(n14928), .Z(n16537) );
  BUF_X1 U12142 ( .A(n14933), .Z(n16513) );
  BUF_X1 U12143 ( .A(n14928), .Z(n16538) );
  BUF_X1 U12144 ( .A(n14933), .Z(n16514) );
  BUF_X1 U12145 ( .A(n14928), .Z(n16539) );
  BUF_X1 U12146 ( .A(n14933), .Z(n16515) );
  BUF_X1 U12147 ( .A(n14928), .Z(n16540) );
  BUF_X1 U12148 ( .A(n14933), .Z(n16516) );
  BUF_X1 U12149 ( .A(n13725), .Z(n16717) );
  BUF_X1 U12150 ( .A(n13725), .Z(n16718) );
  BUF_X1 U12151 ( .A(n13725), .Z(n16719) );
  BUF_X1 U12152 ( .A(n13725), .Z(n16720) );
  BUF_X1 U12153 ( .A(n13725), .Z(n16721) );
  BUF_X1 U12154 ( .A(n14914), .Z(n16583) );
  BUF_X1 U12155 ( .A(n14939), .Z(n16482) );
  BUF_X1 U12156 ( .A(n14914), .Z(n16584) );
  BUF_X1 U12157 ( .A(n14939), .Z(n16483) );
  BUF_X1 U12158 ( .A(n14914), .Z(n16585) );
  BUF_X1 U12159 ( .A(n14939), .Z(n16484) );
  BUF_X1 U12160 ( .A(n14914), .Z(n16586) );
  BUF_X1 U12161 ( .A(n14939), .Z(n16485) );
  BUF_X1 U12162 ( .A(n14914), .Z(n16587) );
  BUF_X1 U12163 ( .A(n14939), .Z(n16486) );
  BUF_X1 U12164 ( .A(n13706), .Z(n16788) );
  BUF_X1 U12165 ( .A(n13731), .Z(n16687) );
  BUF_X1 U12166 ( .A(n13706), .Z(n16789) );
  BUF_X1 U12167 ( .A(n13731), .Z(n16688) );
  BUF_X1 U12168 ( .A(n13706), .Z(n16790) );
  BUF_X1 U12169 ( .A(n13731), .Z(n16689) );
  BUF_X1 U12170 ( .A(n13706), .Z(n16791) );
  BUF_X1 U12171 ( .A(n13731), .Z(n16690) );
  BUF_X1 U12172 ( .A(n13706), .Z(n16792) );
  BUF_X1 U12173 ( .A(n13731), .Z(n16691) );
  BUF_X1 U12174 ( .A(n17580), .Z(n17587) );
  BUF_X1 U12175 ( .A(n17581), .Z(n17588) );
  BUF_X1 U12176 ( .A(n17580), .Z(n17586) );
  BUF_X1 U12177 ( .A(n17580), .Z(n17585) );
  BUF_X1 U12178 ( .A(n17579), .Z(n17584) );
  BUF_X1 U12179 ( .A(n17579), .Z(n17583) );
  BUF_X1 U12180 ( .A(n17579), .Z(n17582) );
  NAND2_X1 U12181 ( .A1(n16082), .A2(n16070), .ZN(n14920) );
  NAND2_X1 U12182 ( .A1(n14874), .A2(n14862), .ZN(n13712) );
  BUF_X1 U12183 ( .A(n14910), .Z(n16605) );
  BUF_X1 U12184 ( .A(n14895), .Z(n16677) );
  BUF_X1 U12185 ( .A(n14900), .Z(n16653) );
  BUF_X1 U12186 ( .A(n14905), .Z(n16629) );
  BUF_X1 U12187 ( .A(n14935), .Z(n16504) );
  BUF_X1 U12188 ( .A(n14930), .Z(n16528) );
  BUF_X1 U12189 ( .A(n13702), .Z(n16810) );
  BUF_X1 U12190 ( .A(n13687), .Z(n16882) );
  BUF_X1 U12191 ( .A(n13692), .Z(n16858) );
  BUF_X1 U12192 ( .A(n13697), .Z(n16834) );
  BUF_X1 U12193 ( .A(n13727), .Z(n16709) );
  BUF_X1 U12194 ( .A(n13722), .Z(n16733) );
  BUF_X1 U12195 ( .A(n14925), .Z(n16548) );
  BUF_X1 U12196 ( .A(n14925), .Z(n16549) );
  BUF_X1 U12197 ( .A(n14925), .Z(n16550) );
  BUF_X1 U12198 ( .A(n14925), .Z(n16551) );
  BUF_X1 U12199 ( .A(n14925), .Z(n16552) );
  BUF_X1 U12200 ( .A(n13717), .Z(n16753) );
  BUF_X1 U12201 ( .A(n13717), .Z(n16754) );
  BUF_X1 U12202 ( .A(n13717), .Z(n16755) );
  BUF_X1 U12203 ( .A(n13717), .Z(n16756) );
  BUF_X1 U12204 ( .A(n13717), .Z(n16757) );
  BUF_X1 U12205 ( .A(n14932), .Z(n16518) );
  BUF_X1 U12206 ( .A(n14909), .Z(n16611) );
  BUF_X1 U12207 ( .A(n14894), .Z(n16683) );
  BUF_X1 U12208 ( .A(n14899), .Z(n16659) );
  BUF_X1 U12209 ( .A(n14904), .Z(n16635) );
  BUF_X1 U12210 ( .A(n14934), .Z(n16510) );
  BUF_X1 U12211 ( .A(n14929), .Z(n16534) );
  BUF_X1 U12212 ( .A(n13701), .Z(n16816) );
  BUF_X1 U12213 ( .A(n13686), .Z(n16888) );
  BUF_X1 U12214 ( .A(n13691), .Z(n16864) );
  BUF_X1 U12215 ( .A(n13696), .Z(n16840) );
  BUF_X1 U12216 ( .A(n13726), .Z(n16715) );
  BUF_X1 U12217 ( .A(n13721), .Z(n16739) );
  BUF_X1 U12218 ( .A(n14924), .Z(n16554) );
  BUF_X1 U12219 ( .A(n14919), .Z(n16577) );
  BUF_X1 U12220 ( .A(n13711), .Z(n16782) );
  BUF_X1 U12221 ( .A(n13716), .Z(n16759) );
  BUF_X1 U12222 ( .A(n17581), .Z(n17589) );
  BUF_X1 U12223 ( .A(n13572), .Z(n17558) );
  OAI21_X1 U12224 ( .B1(n13636), .B2(n13637), .A(n17587), .ZN(n13572) );
  INV_X1 U12225 ( .A(n16890), .ZN(n16906) );
  INV_X1 U12226 ( .A(n16907), .ZN(n16923) );
  INV_X1 U12227 ( .A(n16924), .ZN(n16940) );
  INV_X1 U12228 ( .A(n16941), .ZN(n16957) );
  INV_X1 U12229 ( .A(n16958), .ZN(n16974) );
  INV_X1 U12230 ( .A(n16975), .ZN(n16991) );
  INV_X1 U12231 ( .A(n16992), .ZN(n17008) );
  INV_X1 U12232 ( .A(n17009), .ZN(n17025) );
  INV_X1 U12233 ( .A(n17026), .ZN(n17042) );
  INV_X1 U12234 ( .A(n17043), .ZN(n17059) );
  INV_X1 U12235 ( .A(n17060), .ZN(n17076) );
  INV_X1 U12236 ( .A(n17077), .ZN(n17093) );
  INV_X1 U12237 ( .A(n17094), .ZN(n17110) );
  INV_X1 U12238 ( .A(n17111), .ZN(n17127) );
  INV_X1 U12239 ( .A(n17128), .ZN(n17144) );
  INV_X1 U12240 ( .A(n17145), .ZN(n17161) );
  INV_X1 U12241 ( .A(n17162), .ZN(n17179) );
  INV_X1 U12242 ( .A(n17180), .ZN(n17196) );
  INV_X1 U12243 ( .A(n17197), .ZN(n17213) );
  INV_X1 U12244 ( .A(n17214), .ZN(n17230) );
  INV_X1 U12245 ( .A(n17231), .ZN(n17247) );
  INV_X1 U12246 ( .A(n17248), .ZN(n17264) );
  INV_X1 U12247 ( .A(n17265), .ZN(n17281) );
  INV_X1 U12248 ( .A(n17282), .ZN(n17298) );
  INV_X1 U12249 ( .A(n17299), .ZN(n17317) );
  INV_X1 U12250 ( .A(n17318), .ZN(n17336) );
  INV_X1 U12251 ( .A(n17337), .ZN(n17355) );
  INV_X1 U12252 ( .A(n17356), .ZN(n17374) );
  INV_X1 U12253 ( .A(n17375), .ZN(n17393) );
  INV_X1 U12254 ( .A(n17394), .ZN(n17412) );
  INV_X1 U12255 ( .A(n17413), .ZN(n17431) );
  OAI221_X1 U12256 ( .B1(n13506), .B2(n16530), .C1(n12802), .C2(n16524), .A(
        n16086), .ZN(n16078) );
  AOI22_X1 U12257 ( .A1(n16512), .A2(n12261), .B1(n16547), .B2(n12453), .ZN(
        n16086) );
  OAI221_X1 U12258 ( .B1(n13506), .B2(n16735), .C1(n12802), .C2(n16729), .A(
        n14878), .ZN(n14870) );
  AOI22_X1 U12259 ( .A1(n16723), .A2(n12261), .B1(n16717), .B2(n12453), .ZN(
        n14878) );
  OAI221_X1 U12260 ( .B1(n13505), .B2(n16735), .C1(n12801), .C2(n16729), .A(
        n14846), .ZN(n14841) );
  AOI22_X1 U12261 ( .A1(n16723), .A2(n12260), .B1(n16717), .B2(n12452), .ZN(
        n14846) );
  OAI221_X1 U12262 ( .B1(n13504), .B2(n16735), .C1(n12800), .C2(n16729), .A(
        n14828), .ZN(n14823) );
  AOI22_X1 U12263 ( .A1(n16723), .A2(n12259), .B1(n16717), .B2(n12451), .ZN(
        n14828) );
  OAI221_X1 U12264 ( .B1(n13503), .B2(n16735), .C1(n12799), .C2(n16729), .A(
        n14810), .ZN(n14805) );
  AOI22_X1 U12265 ( .A1(n16723), .A2(n12258), .B1(n16717), .B2(n12450), .ZN(
        n14810) );
  OAI221_X1 U12266 ( .B1(n13502), .B2(n16735), .C1(n12798), .C2(n16729), .A(
        n14792), .ZN(n14787) );
  AOI22_X1 U12267 ( .A1(n16723), .A2(n12257), .B1(n16717), .B2(n12449), .ZN(
        n14792) );
  OAI221_X1 U12268 ( .B1(n13501), .B2(n16735), .C1(n12797), .C2(n16729), .A(
        n14774), .ZN(n14769) );
  AOI22_X1 U12269 ( .A1(n16723), .A2(n12256), .B1(n16717), .B2(n12448), .ZN(
        n14774) );
  OAI221_X1 U12270 ( .B1(n13500), .B2(n16735), .C1(n12796), .C2(n16729), .A(
        n14756), .ZN(n14751) );
  AOI22_X1 U12271 ( .A1(n16723), .A2(n12255), .B1(n16717), .B2(n12447), .ZN(
        n14756) );
  OAI221_X1 U12272 ( .B1(n13499), .B2(n16735), .C1(n12795), .C2(n16729), .A(
        n14738), .ZN(n14733) );
  AOI22_X1 U12273 ( .A1(n16723), .A2(n12254), .B1(n16717), .B2(n12446), .ZN(
        n14738) );
  OAI221_X1 U12274 ( .B1(n13498), .B2(n16735), .C1(n12794), .C2(n16729), .A(
        n14720), .ZN(n14715) );
  AOI22_X1 U12275 ( .A1(n16723), .A2(n12253), .B1(n16717), .B2(n12445), .ZN(
        n14720) );
  OAI221_X1 U12276 ( .B1(n13497), .B2(n16735), .C1(n12793), .C2(n16729), .A(
        n14702), .ZN(n14697) );
  AOI22_X1 U12277 ( .A1(n16723), .A2(n12252), .B1(n16717), .B2(n12444), .ZN(
        n14702) );
  OAI221_X1 U12278 ( .B1(n13496), .B2(n16735), .C1(n12792), .C2(n16729), .A(
        n14684), .ZN(n14679) );
  AOI22_X1 U12279 ( .A1(n16723), .A2(n12251), .B1(n16717), .B2(n12443), .ZN(
        n14684) );
  OAI221_X1 U12280 ( .B1(n13495), .B2(n16735), .C1(n12791), .C2(n16729), .A(
        n14666), .ZN(n14661) );
  AOI22_X1 U12281 ( .A1(n16723), .A2(n12250), .B1(n16717), .B2(n12442), .ZN(
        n14666) );
  OAI221_X1 U12282 ( .B1(n13494), .B2(n16736), .C1(n12790), .C2(n16730), .A(
        n14648), .ZN(n14643) );
  AOI22_X1 U12283 ( .A1(n16724), .A2(n12249), .B1(n16718), .B2(n12441), .ZN(
        n14648) );
  OAI221_X1 U12284 ( .B1(n13493), .B2(n16736), .C1(n12789), .C2(n16730), .A(
        n14630), .ZN(n14625) );
  AOI22_X1 U12285 ( .A1(n16724), .A2(n12248), .B1(n16718), .B2(n12440), .ZN(
        n14630) );
  OAI221_X1 U12286 ( .B1(n13492), .B2(n16736), .C1(n12788), .C2(n16730), .A(
        n14612), .ZN(n14607) );
  AOI22_X1 U12287 ( .A1(n16724), .A2(n12247), .B1(n16718), .B2(n12439), .ZN(
        n14612) );
  OAI221_X1 U12288 ( .B1(n13491), .B2(n16736), .C1(n12787), .C2(n16730), .A(
        n14594), .ZN(n14589) );
  AOI22_X1 U12289 ( .A1(n16724), .A2(n12246), .B1(n16718), .B2(n12438), .ZN(
        n14594) );
  OAI221_X1 U12290 ( .B1(n13490), .B2(n16736), .C1(n12786), .C2(n16730), .A(
        n14576), .ZN(n14571) );
  AOI22_X1 U12291 ( .A1(n16724), .A2(n12245), .B1(n16718), .B2(n12437), .ZN(
        n14576) );
  OAI221_X1 U12292 ( .B1(n13489), .B2(n16736), .C1(n12785), .C2(n16730), .A(
        n14558), .ZN(n14553) );
  AOI22_X1 U12293 ( .A1(n16724), .A2(n12244), .B1(n16718), .B2(n12436), .ZN(
        n14558) );
  OAI221_X1 U12294 ( .B1(n13488), .B2(n16736), .C1(n12784), .C2(n16730), .A(
        n14540), .ZN(n14535) );
  AOI22_X1 U12295 ( .A1(n16724), .A2(n12243), .B1(n16718), .B2(n12435), .ZN(
        n14540) );
  OAI221_X1 U12296 ( .B1(n13487), .B2(n16736), .C1(n12783), .C2(n16730), .A(
        n14522), .ZN(n14517) );
  AOI22_X1 U12297 ( .A1(n16724), .A2(n12242), .B1(n16718), .B2(n12434), .ZN(
        n14522) );
  OAI221_X1 U12298 ( .B1(n13486), .B2(n16736), .C1(n12782), .C2(n16730), .A(
        n14504), .ZN(n14499) );
  AOI22_X1 U12299 ( .A1(n16724), .A2(n12241), .B1(n16718), .B2(n12433), .ZN(
        n14504) );
  OAI221_X1 U12300 ( .B1(n13485), .B2(n16736), .C1(n12781), .C2(n16730), .A(
        n14486), .ZN(n14481) );
  AOI22_X1 U12301 ( .A1(n16724), .A2(n12240), .B1(n16718), .B2(n12432), .ZN(
        n14486) );
  OAI221_X1 U12302 ( .B1(n13484), .B2(n16736), .C1(n12780), .C2(n16730), .A(
        n14468), .ZN(n14463) );
  AOI22_X1 U12303 ( .A1(n16724), .A2(n12239), .B1(n16718), .B2(n12431), .ZN(
        n14468) );
  OAI221_X1 U12304 ( .B1(n13483), .B2(n16736), .C1(n12779), .C2(n16730), .A(
        n14450), .ZN(n14445) );
  AOI22_X1 U12305 ( .A1(n16724), .A2(n12238), .B1(n16718), .B2(n12430), .ZN(
        n14450) );
  OAI221_X1 U12306 ( .B1(n13482), .B2(n16737), .C1(n12778), .C2(n16731), .A(
        n14432), .ZN(n14427) );
  AOI22_X1 U12307 ( .A1(n16725), .A2(n12237), .B1(n16719), .B2(n12429), .ZN(
        n14432) );
  OAI221_X1 U12308 ( .B1(n13481), .B2(n16737), .C1(n12777), .C2(n16731), .A(
        n14414), .ZN(n14409) );
  AOI22_X1 U12309 ( .A1(n16725), .A2(n12236), .B1(n16719), .B2(n12428), .ZN(
        n14414) );
  OAI221_X1 U12310 ( .B1(n13480), .B2(n16737), .C1(n12776), .C2(n16731), .A(
        n14396), .ZN(n14391) );
  AOI22_X1 U12311 ( .A1(n16725), .A2(n12235), .B1(n16719), .B2(n12427), .ZN(
        n14396) );
  OAI221_X1 U12312 ( .B1(n13479), .B2(n16737), .C1(n12775), .C2(n16731), .A(
        n14378), .ZN(n14373) );
  AOI22_X1 U12313 ( .A1(n16725), .A2(n12234), .B1(n16719), .B2(n12426), .ZN(
        n14378) );
  OAI221_X1 U12314 ( .B1(n13478), .B2(n16737), .C1(n12774), .C2(n16731), .A(
        n14360), .ZN(n14355) );
  AOI22_X1 U12315 ( .A1(n16725), .A2(n12233), .B1(n16719), .B2(n12425), .ZN(
        n14360) );
  OAI22_X1 U12316 ( .A1(n17165), .A2(n17437), .B1(n17164), .B2(n12800), .ZN(
        n6030) );
  OAI22_X1 U12317 ( .A1(n17165), .A2(n17439), .B1(n17164), .B2(n12799), .ZN(
        n6031) );
  OAI22_X1 U12318 ( .A1(n17165), .A2(n17441), .B1(n17164), .B2(n12798), .ZN(
        n6032) );
  OAI22_X1 U12319 ( .A1(n17166), .A2(n17443), .B1(n17164), .B2(n12797), .ZN(
        n6033) );
  OAI22_X1 U12320 ( .A1(n17166), .A2(n17445), .B1(n17164), .B2(n12796), .ZN(
        n6034) );
  OAI22_X1 U12321 ( .A1(n17166), .A2(n17447), .B1(n17164), .B2(n12795), .ZN(
        n6035) );
  OAI22_X1 U12322 ( .A1(n17166), .A2(n17449), .B1(n17164), .B2(n12794), .ZN(
        n6036) );
  OAI22_X1 U12323 ( .A1(n17166), .A2(n17451), .B1(n17164), .B2(n12793), .ZN(
        n6037) );
  OAI22_X1 U12324 ( .A1(n17167), .A2(n17453), .B1(n17164), .B2(n12792), .ZN(
        n6038) );
  OAI22_X1 U12325 ( .A1(n17167), .A2(n17455), .B1(n17164), .B2(n12791), .ZN(
        n6039) );
  OAI22_X1 U12326 ( .A1(n17167), .A2(n17457), .B1(n17164), .B2(n12790), .ZN(
        n6040) );
  OAI22_X1 U12327 ( .A1(n17167), .A2(n17459), .B1(n17164), .B2(n12789), .ZN(
        n6041) );
  OAI22_X1 U12328 ( .A1(n17167), .A2(n17461), .B1(n17164), .B2(n12788), .ZN(
        n6042) );
  OAI22_X1 U12329 ( .A1(n17168), .A2(n17463), .B1(n17164), .B2(n12787), .ZN(
        n6043) );
  OAI22_X1 U12330 ( .A1(n17168), .A2(n17465), .B1(n17163), .B2(n12786), .ZN(
        n6044) );
  OAI22_X1 U12331 ( .A1(n17168), .A2(n17467), .B1(n17162), .B2(n12785), .ZN(
        n6045) );
  OAI22_X1 U12332 ( .A1(n17168), .A2(n17469), .B1(n17164), .B2(n12784), .ZN(
        n6046) );
  OAI22_X1 U12333 ( .A1(n17168), .A2(n17471), .B1(n17163), .B2(n12783), .ZN(
        n6047) );
  OAI22_X1 U12334 ( .A1(n17169), .A2(n17473), .B1(n17162), .B2(n12782), .ZN(
        n6048) );
  OAI22_X1 U12335 ( .A1(n17169), .A2(n17475), .B1(n17164), .B2(n12781), .ZN(
        n6049) );
  OAI22_X1 U12336 ( .A1(n17169), .A2(n17477), .B1(n17163), .B2(n12780), .ZN(
        n6050) );
  OAI22_X1 U12337 ( .A1(n17169), .A2(n17479), .B1(n17162), .B2(n12779), .ZN(
        n6051) );
  OAI22_X1 U12338 ( .A1(n17169), .A2(n17481), .B1(n17164), .B2(n12778), .ZN(
        n6052) );
  OAI22_X1 U12339 ( .A1(n17170), .A2(n17483), .B1(n17163), .B2(n12777), .ZN(
        n6053) );
  OAI22_X1 U12340 ( .A1(n17170), .A2(n17485), .B1(n17162), .B2(n12776), .ZN(
        n6054) );
  OAI22_X1 U12341 ( .A1(n17170), .A2(n17487), .B1(n17164), .B2(n12775), .ZN(
        n6055) );
  OAI22_X1 U12342 ( .A1(n17170), .A2(n17489), .B1(n17163), .B2(n12774), .ZN(
        n6056) );
  OAI22_X1 U12343 ( .A1(n16893), .A2(n17432), .B1(n16891), .B2(n13570), .ZN(
        n5004) );
  OAI22_X1 U12344 ( .A1(n16893), .A2(n17434), .B1(n16891), .B2(n13569), .ZN(
        n5005) );
  OAI22_X1 U12345 ( .A1(n16893), .A2(n17436), .B1(n16891), .B2(n13568), .ZN(
        n5006) );
  OAI22_X1 U12346 ( .A1(n16893), .A2(n17438), .B1(n16891), .B2(n13567), .ZN(
        n5007) );
  OAI22_X1 U12347 ( .A1(n16893), .A2(n17440), .B1(n16891), .B2(n13566), .ZN(
        n5008) );
  OAI22_X1 U12348 ( .A1(n16894), .A2(n17442), .B1(n16891), .B2(n13565), .ZN(
        n5009) );
  OAI22_X1 U12349 ( .A1(n16894), .A2(n17444), .B1(n16891), .B2(n13564), .ZN(
        n5010) );
  OAI22_X1 U12350 ( .A1(n16894), .A2(n17446), .B1(n16891), .B2(n13563), .ZN(
        n5011) );
  OAI22_X1 U12351 ( .A1(n16894), .A2(n17448), .B1(n16891), .B2(n13562), .ZN(
        n5012) );
  OAI22_X1 U12352 ( .A1(n16894), .A2(n17450), .B1(n16891), .B2(n13561), .ZN(
        n5013) );
  OAI22_X1 U12353 ( .A1(n16895), .A2(n17452), .B1(n16891), .B2(n13560), .ZN(
        n5014) );
  OAI22_X1 U12354 ( .A1(n16895), .A2(n17454), .B1(n16891), .B2(n13559), .ZN(
        n5015) );
  OAI22_X1 U12355 ( .A1(n16895), .A2(n17456), .B1(n16892), .B2(n13558), .ZN(
        n5016) );
  OAI22_X1 U12356 ( .A1(n16895), .A2(n17458), .B1(n16892), .B2(n13557), .ZN(
        n5017) );
  OAI22_X1 U12357 ( .A1(n16895), .A2(n17460), .B1(n16892), .B2(n13556), .ZN(
        n5018) );
  OAI22_X1 U12358 ( .A1(n16896), .A2(n17462), .B1(n16892), .B2(n13555), .ZN(
        n5019) );
  OAI22_X1 U12359 ( .A1(n16896), .A2(n17464), .B1(n16892), .B2(n13554), .ZN(
        n5020) );
  OAI22_X1 U12360 ( .A1(n16896), .A2(n17466), .B1(n16892), .B2(n13553), .ZN(
        n5021) );
  OAI22_X1 U12361 ( .A1(n16896), .A2(n17468), .B1(n16892), .B2(n13552), .ZN(
        n5022) );
  OAI22_X1 U12362 ( .A1(n16896), .A2(n17470), .B1(n16892), .B2(n13551), .ZN(
        n5023) );
  OAI22_X1 U12363 ( .A1(n16897), .A2(n17472), .B1(n16892), .B2(n13550), .ZN(
        n5024) );
  OAI22_X1 U12364 ( .A1(n16897), .A2(n17474), .B1(n16892), .B2(n13549), .ZN(
        n5025) );
  OAI22_X1 U12365 ( .A1(n16897), .A2(n17476), .B1(n16892), .B2(n13548), .ZN(
        n5026) );
  OAI22_X1 U12366 ( .A1(n16897), .A2(n17478), .B1(n16892), .B2(n13547), .ZN(
        n5027) );
  OAI22_X1 U12367 ( .A1(n16910), .A2(n17432), .B1(n16908), .B2(n13506), .ZN(
        n5068) );
  OAI22_X1 U12368 ( .A1(n16910), .A2(n17434), .B1(n16908), .B2(n13505), .ZN(
        n5069) );
  OAI22_X1 U12369 ( .A1(n16910), .A2(n17436), .B1(n16908), .B2(n13504), .ZN(
        n5070) );
  OAI22_X1 U12370 ( .A1(n16910), .A2(n17438), .B1(n16908), .B2(n13503), .ZN(
        n5071) );
  OAI22_X1 U12371 ( .A1(n16910), .A2(n17440), .B1(n16908), .B2(n13502), .ZN(
        n5072) );
  OAI22_X1 U12372 ( .A1(n16911), .A2(n17442), .B1(n16908), .B2(n13501), .ZN(
        n5073) );
  OAI22_X1 U12373 ( .A1(n16911), .A2(n17444), .B1(n16908), .B2(n13500), .ZN(
        n5074) );
  OAI22_X1 U12374 ( .A1(n16911), .A2(n17446), .B1(n16908), .B2(n13499), .ZN(
        n5075) );
  OAI22_X1 U12375 ( .A1(n16911), .A2(n17448), .B1(n16908), .B2(n13498), .ZN(
        n5076) );
  OAI22_X1 U12376 ( .A1(n16911), .A2(n17450), .B1(n16908), .B2(n13497), .ZN(
        n5077) );
  OAI22_X1 U12377 ( .A1(n16912), .A2(n17452), .B1(n16908), .B2(n13496), .ZN(
        n5078) );
  OAI22_X1 U12378 ( .A1(n16912), .A2(n17454), .B1(n16908), .B2(n13495), .ZN(
        n5079) );
  OAI22_X1 U12379 ( .A1(n16912), .A2(n17456), .B1(n16909), .B2(n13494), .ZN(
        n5080) );
  OAI22_X1 U12380 ( .A1(n16912), .A2(n17458), .B1(n16909), .B2(n13493), .ZN(
        n5081) );
  OAI22_X1 U12381 ( .A1(n16912), .A2(n17460), .B1(n16909), .B2(n13492), .ZN(
        n5082) );
  OAI22_X1 U12382 ( .A1(n16913), .A2(n17462), .B1(n16909), .B2(n13491), .ZN(
        n5083) );
  OAI22_X1 U12383 ( .A1(n16913), .A2(n17464), .B1(n16909), .B2(n13490), .ZN(
        n5084) );
  OAI22_X1 U12384 ( .A1(n16913), .A2(n17466), .B1(n16909), .B2(n13489), .ZN(
        n5085) );
  OAI22_X1 U12385 ( .A1(n16913), .A2(n17468), .B1(n16909), .B2(n13488), .ZN(
        n5086) );
  OAI22_X1 U12386 ( .A1(n16913), .A2(n17470), .B1(n16909), .B2(n13487), .ZN(
        n5087) );
  OAI22_X1 U12387 ( .A1(n16914), .A2(n17472), .B1(n16909), .B2(n13486), .ZN(
        n5088) );
  OAI22_X1 U12388 ( .A1(n16914), .A2(n17474), .B1(n16909), .B2(n13485), .ZN(
        n5089) );
  OAI22_X1 U12389 ( .A1(n16914), .A2(n17476), .B1(n16909), .B2(n13484), .ZN(
        n5090) );
  OAI22_X1 U12390 ( .A1(n16914), .A2(n17478), .B1(n16909), .B2(n13483), .ZN(
        n5091) );
  OAI22_X1 U12391 ( .A1(n17063), .A2(n17432), .B1(n17061), .B2(n13058), .ZN(
        n5644) );
  OAI22_X1 U12392 ( .A1(n17063), .A2(n17434), .B1(n17061), .B2(n13057), .ZN(
        n5645) );
  OAI22_X1 U12393 ( .A1(n17063), .A2(n17436), .B1(n17061), .B2(n13056), .ZN(
        n5646) );
  OAI22_X1 U12394 ( .A1(n17063), .A2(n17438), .B1(n17061), .B2(n13055), .ZN(
        n5647) );
  OAI22_X1 U12395 ( .A1(n17063), .A2(n17440), .B1(n17061), .B2(n13054), .ZN(
        n5648) );
  OAI22_X1 U12396 ( .A1(n17064), .A2(n17442), .B1(n17061), .B2(n13053), .ZN(
        n5649) );
  OAI22_X1 U12397 ( .A1(n17064), .A2(n17444), .B1(n17061), .B2(n13052), .ZN(
        n5650) );
  OAI22_X1 U12398 ( .A1(n17064), .A2(n17446), .B1(n17061), .B2(n13051), .ZN(
        n5651) );
  OAI22_X1 U12399 ( .A1(n17064), .A2(n17448), .B1(n17061), .B2(n13050), .ZN(
        n5652) );
  OAI22_X1 U12400 ( .A1(n17064), .A2(n17450), .B1(n17061), .B2(n13049), .ZN(
        n5653) );
  OAI22_X1 U12401 ( .A1(n17065), .A2(n17452), .B1(n17061), .B2(n13048), .ZN(
        n5654) );
  OAI22_X1 U12402 ( .A1(n17065), .A2(n17454), .B1(n17061), .B2(n13047), .ZN(
        n5655) );
  OAI22_X1 U12403 ( .A1(n17065), .A2(n17456), .B1(n17062), .B2(n13046), .ZN(
        n5656) );
  OAI22_X1 U12404 ( .A1(n17065), .A2(n17458), .B1(n17062), .B2(n13045), .ZN(
        n5657) );
  OAI22_X1 U12405 ( .A1(n17065), .A2(n17460), .B1(n17062), .B2(n13044), .ZN(
        n5658) );
  OAI22_X1 U12406 ( .A1(n17066), .A2(n17462), .B1(n17062), .B2(n13043), .ZN(
        n5659) );
  OAI22_X1 U12407 ( .A1(n17066), .A2(n17464), .B1(n17062), .B2(n13042), .ZN(
        n5660) );
  OAI22_X1 U12408 ( .A1(n17066), .A2(n17466), .B1(n17062), .B2(n13041), .ZN(
        n5661) );
  OAI22_X1 U12409 ( .A1(n17066), .A2(n17468), .B1(n17062), .B2(n13040), .ZN(
        n5662) );
  OAI22_X1 U12410 ( .A1(n17066), .A2(n17470), .B1(n17062), .B2(n13039), .ZN(
        n5663) );
  OAI22_X1 U12411 ( .A1(n17067), .A2(n17472), .B1(n17062), .B2(n13038), .ZN(
        n5664) );
  OAI22_X1 U12412 ( .A1(n17067), .A2(n17474), .B1(n17062), .B2(n13037), .ZN(
        n5665) );
  OAI22_X1 U12413 ( .A1(n17067), .A2(n17476), .B1(n17062), .B2(n13036), .ZN(
        n5666) );
  OAI22_X1 U12414 ( .A1(n17067), .A2(n17478), .B1(n17062), .B2(n13035), .ZN(
        n5667) );
  OAI22_X1 U12415 ( .A1(n17217), .A2(n17433), .B1(n17215), .B2(n12773), .ZN(
        n6220) );
  OAI22_X1 U12416 ( .A1(n17217), .A2(n17435), .B1(n17215), .B2(n12772), .ZN(
        n6221) );
  OAI22_X1 U12417 ( .A1(n17217), .A2(n17437), .B1(n17215), .B2(n12771), .ZN(
        n6222) );
  OAI22_X1 U12418 ( .A1(n17217), .A2(n17439), .B1(n17215), .B2(n12770), .ZN(
        n6223) );
  OAI22_X1 U12419 ( .A1(n17217), .A2(n17441), .B1(n17215), .B2(n12769), .ZN(
        n6224) );
  OAI22_X1 U12420 ( .A1(n17218), .A2(n17443), .B1(n17215), .B2(n12768), .ZN(
        n6225) );
  OAI22_X1 U12421 ( .A1(n17218), .A2(n17445), .B1(n17215), .B2(n12767), .ZN(
        n6226) );
  OAI22_X1 U12422 ( .A1(n17218), .A2(n17447), .B1(n17215), .B2(n12766), .ZN(
        n6227) );
  OAI22_X1 U12423 ( .A1(n17218), .A2(n17449), .B1(n17215), .B2(n12765), .ZN(
        n6228) );
  OAI22_X1 U12424 ( .A1(n17218), .A2(n17451), .B1(n17215), .B2(n12764), .ZN(
        n6229) );
  OAI22_X1 U12425 ( .A1(n17219), .A2(n17453), .B1(n17215), .B2(n12763), .ZN(
        n6230) );
  OAI22_X1 U12426 ( .A1(n17219), .A2(n17455), .B1(n17215), .B2(n12762), .ZN(
        n6231) );
  OAI22_X1 U12427 ( .A1(n17219), .A2(n17457), .B1(n17216), .B2(n12761), .ZN(
        n6232) );
  OAI22_X1 U12428 ( .A1(n17219), .A2(n17459), .B1(n17216), .B2(n12760), .ZN(
        n6233) );
  OAI22_X1 U12429 ( .A1(n17219), .A2(n17461), .B1(n17216), .B2(n12759), .ZN(
        n6234) );
  OAI22_X1 U12430 ( .A1(n17220), .A2(n17463), .B1(n17216), .B2(n12758), .ZN(
        n6235) );
  OAI22_X1 U12431 ( .A1(n17220), .A2(n17465), .B1(n17216), .B2(n12757), .ZN(
        n6236) );
  OAI22_X1 U12432 ( .A1(n17220), .A2(n17467), .B1(n17216), .B2(n12756), .ZN(
        n6237) );
  OAI22_X1 U12433 ( .A1(n17220), .A2(n17469), .B1(n17216), .B2(n12755), .ZN(
        n6238) );
  OAI22_X1 U12434 ( .A1(n17220), .A2(n17471), .B1(n17216), .B2(n12754), .ZN(
        n6239) );
  OAI22_X1 U12435 ( .A1(n17221), .A2(n17473), .B1(n17216), .B2(n12753), .ZN(
        n6240) );
  OAI22_X1 U12436 ( .A1(n17221), .A2(n17475), .B1(n17216), .B2(n12752), .ZN(
        n6241) );
  OAI22_X1 U12437 ( .A1(n17221), .A2(n17477), .B1(n17216), .B2(n12751), .ZN(
        n6242) );
  OAI22_X1 U12438 ( .A1(n17221), .A2(n17479), .B1(n17216), .B2(n12750), .ZN(
        n6243) );
  OAI22_X1 U12439 ( .A1(n17251), .A2(n17433), .B1(n17249), .B2(n12645), .ZN(
        n6348) );
  OAI22_X1 U12440 ( .A1(n17251), .A2(n17435), .B1(n17249), .B2(n12644), .ZN(
        n6349) );
  OAI22_X1 U12441 ( .A1(n17251), .A2(n17437), .B1(n17249), .B2(n12643), .ZN(
        n6350) );
  OAI22_X1 U12442 ( .A1(n17251), .A2(n17439), .B1(n17249), .B2(n12642), .ZN(
        n6351) );
  OAI22_X1 U12443 ( .A1(n17251), .A2(n17441), .B1(n17249), .B2(n12641), .ZN(
        n6352) );
  OAI22_X1 U12444 ( .A1(n17252), .A2(n17443), .B1(n17249), .B2(n12640), .ZN(
        n6353) );
  OAI22_X1 U12445 ( .A1(n17252), .A2(n17445), .B1(n17249), .B2(n12639), .ZN(
        n6354) );
  OAI22_X1 U12446 ( .A1(n17252), .A2(n17447), .B1(n17249), .B2(n12638), .ZN(
        n6355) );
  OAI22_X1 U12447 ( .A1(n17252), .A2(n17449), .B1(n17249), .B2(n12637), .ZN(
        n6356) );
  OAI22_X1 U12448 ( .A1(n17252), .A2(n17451), .B1(n17249), .B2(n12636), .ZN(
        n6357) );
  OAI22_X1 U12449 ( .A1(n17253), .A2(n17453), .B1(n17249), .B2(n12635), .ZN(
        n6358) );
  OAI22_X1 U12450 ( .A1(n17253), .A2(n17455), .B1(n17249), .B2(n12634), .ZN(
        n6359) );
  OAI22_X1 U12451 ( .A1(n17253), .A2(n17457), .B1(n17250), .B2(n12633), .ZN(
        n6360) );
  OAI22_X1 U12452 ( .A1(n17253), .A2(n17459), .B1(n17250), .B2(n12632), .ZN(
        n6361) );
  OAI22_X1 U12453 ( .A1(n17253), .A2(n17461), .B1(n17250), .B2(n12631), .ZN(
        n6362) );
  OAI22_X1 U12454 ( .A1(n17254), .A2(n17463), .B1(n17250), .B2(n12630), .ZN(
        n6363) );
  OAI22_X1 U12455 ( .A1(n17254), .A2(n17465), .B1(n17250), .B2(n12629), .ZN(
        n6364) );
  OAI22_X1 U12456 ( .A1(n17254), .A2(n17467), .B1(n17250), .B2(n12628), .ZN(
        n6365) );
  OAI22_X1 U12457 ( .A1(n17254), .A2(n17469), .B1(n17250), .B2(n12627), .ZN(
        n6366) );
  OAI22_X1 U12458 ( .A1(n17254), .A2(n17471), .B1(n17250), .B2(n12626), .ZN(
        n6367) );
  OAI22_X1 U12459 ( .A1(n17255), .A2(n17473), .B1(n17250), .B2(n12625), .ZN(
        n6368) );
  OAI22_X1 U12460 ( .A1(n17255), .A2(n17475), .B1(n17250), .B2(n12624), .ZN(
        n6369) );
  OAI22_X1 U12461 ( .A1(n17255), .A2(n17477), .B1(n17250), .B2(n12623), .ZN(
        n6370) );
  OAI22_X1 U12462 ( .A1(n17255), .A2(n17479), .B1(n17250), .B2(n12622), .ZN(
        n6371) );
  AOI22_X1 U12463 ( .A1(n16536), .A2(n12325), .B1(n16523), .B2(n16479), .ZN(
        n16084) );
  AOI22_X1 U12464 ( .A1(n16523), .A2(n16420), .B1(n16512), .B2(n12260), .ZN(
        n16054) );
  AOI22_X1 U12465 ( .A1(n16523), .A2(n16421), .B1(n16512), .B2(n12259), .ZN(
        n16036) );
  AOI22_X1 U12466 ( .A1(n16523), .A2(n16422), .B1(n16512), .B2(n12258), .ZN(
        n16018) );
  AOI22_X1 U12467 ( .A1(n16522), .A2(n16423), .B1(n16512), .B2(n12257), .ZN(
        n16000) );
  AOI22_X1 U12468 ( .A1(n16522), .A2(n16424), .B1(n16512), .B2(n12256), .ZN(
        n15982) );
  AOI22_X1 U12469 ( .A1(n16522), .A2(n16425), .B1(n16512), .B2(n12255), .ZN(
        n15964) );
  AOI22_X1 U12470 ( .A1(n16522), .A2(n16426), .B1(n16512), .B2(n12254), .ZN(
        n15946) );
  AOI22_X1 U12471 ( .A1(n16522), .A2(n16427), .B1(n16512), .B2(n12253), .ZN(
        n15928) );
  AOI22_X1 U12472 ( .A1(n16522), .A2(n16428), .B1(n16512), .B2(n12252), .ZN(
        n15910) );
  AOI22_X1 U12473 ( .A1(n16522), .A2(n16429), .B1(n16512), .B2(n12251), .ZN(
        n15892) );
  AOI22_X1 U12474 ( .A1(n16522), .A2(n16430), .B1(n16512), .B2(n12250), .ZN(
        n15874) );
  AOI22_X1 U12475 ( .A1(n16522), .A2(n16431), .B1(n16513), .B2(n12249), .ZN(
        n15856) );
  AOI22_X1 U12476 ( .A1(n16522), .A2(n16432), .B1(n16513), .B2(n12248), .ZN(
        n15838) );
  AOI22_X1 U12477 ( .A1(n16522), .A2(n16433), .B1(n16513), .B2(n12247), .ZN(
        n15820) );
  AOI22_X1 U12478 ( .A1(n16522), .A2(n16434), .B1(n16513), .B2(n12246), .ZN(
        n15802) );
  AOI22_X1 U12479 ( .A1(n16521), .A2(n16435), .B1(n16513), .B2(n12245), .ZN(
        n15784) );
  AOI22_X1 U12480 ( .A1(n16521), .A2(n16436), .B1(n16513), .B2(n12244), .ZN(
        n15766) );
  AOI22_X1 U12481 ( .A1(n16521), .A2(n16437), .B1(n16513), .B2(n12243), .ZN(
        n15748) );
  AOI22_X1 U12482 ( .A1(n16521), .A2(n16438), .B1(n16513), .B2(n12242), .ZN(
        n15730) );
  AOI22_X1 U12483 ( .A1(n16521), .A2(n16439), .B1(n16513), .B2(n12241), .ZN(
        n15712) );
  AOI22_X1 U12484 ( .A1(n16521), .A2(n16440), .B1(n16513), .B2(n12240), .ZN(
        n15694) );
  AOI22_X1 U12485 ( .A1(n16521), .A2(n16441), .B1(n16513), .B2(n12239), .ZN(
        n15676) );
  AOI22_X1 U12486 ( .A1(n16521), .A2(n16442), .B1(n16513), .B2(n12238), .ZN(
        n15658) );
  AOI22_X1 U12487 ( .A1(n16521), .A2(n16443), .B1(n16514), .B2(n12237), .ZN(
        n15640) );
  AOI22_X1 U12488 ( .A1(n16521), .A2(n16444), .B1(n16514), .B2(n12236), .ZN(
        n15622) );
  AOI22_X1 U12489 ( .A1(n16521), .A2(n16445), .B1(n16514), .B2(n12235), .ZN(
        n15604) );
  AOI22_X1 U12490 ( .A1(n16521), .A2(n16446), .B1(n16514), .B2(n12234), .ZN(
        n15586) );
  AOI22_X1 U12491 ( .A1(n16520), .A2(n16447), .B1(n16514), .B2(n12233), .ZN(
        n15568) );
  AOI22_X1 U12492 ( .A1(n16520), .A2(n16448), .B1(n16514), .B2(n12232), .ZN(
        n15550) );
  AOI22_X1 U12493 ( .A1(n16520), .A2(n16449), .B1(n16514), .B2(n12231), .ZN(
        n15532) );
  AOI22_X1 U12494 ( .A1(n16520), .A2(n16450), .B1(n16514), .B2(n12230), .ZN(
        n15514) );
  AOI22_X1 U12495 ( .A1(n16520), .A2(n16451), .B1(n16514), .B2(n12229), .ZN(
        n15496) );
  AOI22_X1 U12496 ( .A1(n16520), .A2(n16452), .B1(n16514), .B2(n12228), .ZN(
        n15478) );
  AOI22_X1 U12497 ( .A1(n16520), .A2(n16453), .B1(n16514), .B2(n12227), .ZN(
        n15460) );
  AOI22_X1 U12498 ( .A1(n16520), .A2(n16454), .B1(n16514), .B2(n12226), .ZN(
        n15442) );
  AOI22_X1 U12499 ( .A1(n16520), .A2(n16455), .B1(n16515), .B2(n12225), .ZN(
        n15424) );
  AOI22_X1 U12500 ( .A1(n16520), .A2(n16456), .B1(n16515), .B2(n12224), .ZN(
        n15406) );
  AOI22_X1 U12501 ( .A1(n16520), .A2(n16457), .B1(n16515), .B2(n12223), .ZN(
        n15388) );
  AOI22_X1 U12502 ( .A1(n16520), .A2(n16458), .B1(n16515), .B2(n12222), .ZN(
        n15370) );
  AOI22_X1 U12503 ( .A1(n16519), .A2(n16459), .B1(n16515), .B2(n12221), .ZN(
        n15352) );
  AOI22_X1 U12504 ( .A1(n16519), .A2(n16460), .B1(n16515), .B2(n12220), .ZN(
        n15334) );
  AOI22_X1 U12505 ( .A1(n16519), .A2(n16461), .B1(n16515), .B2(n12219), .ZN(
        n15316) );
  AOI22_X1 U12506 ( .A1(n16519), .A2(n16462), .B1(n16515), .B2(n12218), .ZN(
        n15298) );
  AOI22_X1 U12507 ( .A1(n16519), .A2(n16463), .B1(n16515), .B2(n12217), .ZN(
        n15280) );
  AOI22_X1 U12508 ( .A1(n16519), .A2(n16464), .B1(n16515), .B2(n12216), .ZN(
        n15262) );
  AOI22_X1 U12509 ( .A1(n16519), .A2(n16465), .B1(n16515), .B2(n12215), .ZN(
        n15244) );
  AOI22_X1 U12510 ( .A1(n16519), .A2(n16466), .B1(n16515), .B2(n12214), .ZN(
        n15226) );
  AOI22_X1 U12511 ( .A1(n16519), .A2(n16467), .B1(n16516), .B2(n12213), .ZN(
        n15208) );
  AOI22_X1 U12512 ( .A1(n16519), .A2(n16468), .B1(n16516), .B2(n12212), .ZN(
        n15190) );
  AOI22_X1 U12513 ( .A1(n16519), .A2(n16469), .B1(n16516), .B2(n12211), .ZN(
        n15172) );
  AOI22_X1 U12514 ( .A1(n16519), .A2(n16470), .B1(n16516), .B2(n12210), .ZN(
        n15154) );
  AOI22_X1 U12515 ( .A1(n16518), .A2(n16471), .B1(n16516), .B2(n12209), .ZN(
        n15136) );
  AOI22_X1 U12516 ( .A1(n16518), .A2(n16472), .B1(n16516), .B2(n12208), .ZN(
        n15118) );
  AOI22_X1 U12517 ( .A1(n16518), .A2(n16473), .B1(n16516), .B2(n12207), .ZN(
        n15100) );
  AOI22_X1 U12518 ( .A1(n16518), .A2(n16474), .B1(n16516), .B2(n12206), .ZN(
        n15082) );
  AOI22_X1 U12519 ( .A1(n16518), .A2(n16475), .B1(n16516), .B2(n12205), .ZN(
        n15064) );
  AOI22_X1 U12520 ( .A1(n16518), .A2(n16476), .B1(n16516), .B2(n12204), .ZN(
        n15046) );
  AOI22_X1 U12521 ( .A1(n16518), .A2(n16477), .B1(n16516), .B2(n12203), .ZN(
        n15028) );
  AOI22_X1 U12522 ( .A1(n16518), .A2(n16478), .B1(n16516), .B2(n12202), .ZN(
        n15010) );
  AOI22_X1 U12523 ( .A1(n16518), .A2(n16416), .B1(n16517), .B2(n12201), .ZN(
        n14992) );
  AOI22_X1 U12524 ( .A1(n16518), .A2(n16417), .B1(n16517), .B2(n12200), .ZN(
        n14974) );
  AOI22_X1 U12525 ( .A1(n16518), .A2(n16418), .B1(n16517), .B2(n12199), .ZN(
        n14956) );
  AOI22_X1 U12526 ( .A1(n16518), .A2(n16419), .B1(n16517), .B2(n12198), .ZN(
        n14931) );
  AOI22_X1 U12527 ( .A1(n16747), .A2(n12325), .B1(n16741), .B2(n16479), .ZN(
        n14876) );
  AOI22_X1 U12528 ( .A1(n16747), .A2(n12324), .B1(n16741), .B2(n16420), .ZN(
        n14845) );
  AOI22_X1 U12529 ( .A1(n16747), .A2(n12323), .B1(n16741), .B2(n16421), .ZN(
        n14827) );
  AOI22_X1 U12530 ( .A1(n16747), .A2(n12322), .B1(n16741), .B2(n16422), .ZN(
        n14809) );
  AOI22_X1 U12531 ( .A1(n16747), .A2(n12321), .B1(n16741), .B2(n16423), .ZN(
        n14791) );
  AOI22_X1 U12532 ( .A1(n16747), .A2(n12320), .B1(n16741), .B2(n16424), .ZN(
        n14773) );
  AOI22_X1 U12533 ( .A1(n16747), .A2(n12319), .B1(n16741), .B2(n16425), .ZN(
        n14755) );
  AOI22_X1 U12534 ( .A1(n16747), .A2(n12318), .B1(n16741), .B2(n16426), .ZN(
        n14737) );
  AOI22_X1 U12535 ( .A1(n16747), .A2(n12317), .B1(n16741), .B2(n16427), .ZN(
        n14719) );
  AOI22_X1 U12536 ( .A1(n16747), .A2(n12316), .B1(n16741), .B2(n16428), .ZN(
        n14701) );
  AOI22_X1 U12537 ( .A1(n16747), .A2(n12315), .B1(n16741), .B2(n16429), .ZN(
        n14683) );
  AOI22_X1 U12538 ( .A1(n16747), .A2(n12314), .B1(n16741), .B2(n16430), .ZN(
        n14665) );
  AOI22_X1 U12539 ( .A1(n16748), .A2(n12313), .B1(n16742), .B2(n16431), .ZN(
        n14647) );
  AOI22_X1 U12540 ( .A1(n16748), .A2(n12312), .B1(n16742), .B2(n16432), .ZN(
        n14629) );
  AOI22_X1 U12541 ( .A1(n16748), .A2(n12311), .B1(n16742), .B2(n16433), .ZN(
        n14611) );
  AOI22_X1 U12542 ( .A1(n16748), .A2(n12310), .B1(n16742), .B2(n16434), .ZN(
        n14593) );
  AOI22_X1 U12543 ( .A1(n16748), .A2(n12309), .B1(n16742), .B2(n16435), .ZN(
        n14575) );
  AOI22_X1 U12544 ( .A1(n16748), .A2(n12308), .B1(n16742), .B2(n16436), .ZN(
        n14557) );
  AOI22_X1 U12545 ( .A1(n16748), .A2(n12307), .B1(n16742), .B2(n16437), .ZN(
        n14539) );
  AOI22_X1 U12546 ( .A1(n16748), .A2(n12306), .B1(n16742), .B2(n16438), .ZN(
        n14521) );
  AOI22_X1 U12547 ( .A1(n16748), .A2(n12305), .B1(n16742), .B2(n16439), .ZN(
        n14503) );
  AOI22_X1 U12548 ( .A1(n16748), .A2(n12304), .B1(n16742), .B2(n16440), .ZN(
        n14485) );
  AOI22_X1 U12549 ( .A1(n16748), .A2(n12303), .B1(n16742), .B2(n16441), .ZN(
        n14467) );
  AOI22_X1 U12550 ( .A1(n16748), .A2(n12302), .B1(n16742), .B2(n16442), .ZN(
        n14449) );
  AOI22_X1 U12551 ( .A1(n16749), .A2(n12301), .B1(n16743), .B2(n16443), .ZN(
        n14431) );
  AOI22_X1 U12552 ( .A1(n16749), .A2(n12300), .B1(n16743), .B2(n16444), .ZN(
        n14413) );
  AOI22_X1 U12553 ( .A1(n16749), .A2(n12299), .B1(n16743), .B2(n16445), .ZN(
        n14395) );
  AOI22_X1 U12554 ( .A1(n16749), .A2(n12298), .B1(n16743), .B2(n16446), .ZN(
        n14377) );
  AOI22_X1 U12555 ( .A1(n16749), .A2(n12297), .B1(n16743), .B2(n16447), .ZN(
        n14359) );
  AOI22_X1 U12556 ( .A1(n16749), .A2(n12296), .B1(n16743), .B2(n16448), .ZN(
        n14341) );
  AOI22_X1 U12557 ( .A1(n16749), .A2(n12295), .B1(n16743), .B2(n16449), .ZN(
        n14323) );
  AOI22_X1 U12558 ( .A1(n16749), .A2(n12294), .B1(n16743), .B2(n16450), .ZN(
        n14305) );
  AOI22_X1 U12559 ( .A1(n16749), .A2(n12293), .B1(n16743), .B2(n16451), .ZN(
        n14287) );
  AOI22_X1 U12560 ( .A1(n16749), .A2(n12292), .B1(n16743), .B2(n16452), .ZN(
        n14269) );
  AOI22_X1 U12561 ( .A1(n16749), .A2(n12291), .B1(n16743), .B2(n16453), .ZN(
        n14251) );
  AOI22_X1 U12562 ( .A1(n16749), .A2(n12290), .B1(n16743), .B2(n16454), .ZN(
        n14233) );
  AOI22_X1 U12563 ( .A1(n16750), .A2(n12289), .B1(n16744), .B2(n16455), .ZN(
        n14215) );
  AOI22_X1 U12564 ( .A1(n16750), .A2(n12288), .B1(n16744), .B2(n16456), .ZN(
        n14197) );
  AOI22_X1 U12565 ( .A1(n16750), .A2(n12287), .B1(n16744), .B2(n16457), .ZN(
        n14179) );
  AOI22_X1 U12566 ( .A1(n16750), .A2(n12286), .B1(n16744), .B2(n16458), .ZN(
        n14161) );
  AOI22_X1 U12567 ( .A1(n16750), .A2(n12285), .B1(n16744), .B2(n16459), .ZN(
        n14143) );
  AOI22_X1 U12568 ( .A1(n16750), .A2(n12284), .B1(n16744), .B2(n16460), .ZN(
        n14125) );
  AOI22_X1 U12569 ( .A1(n16750), .A2(n12283), .B1(n16744), .B2(n16461), .ZN(
        n14107) );
  AOI22_X1 U12570 ( .A1(n16750), .A2(n12282), .B1(n16744), .B2(n16462), .ZN(
        n14089) );
  AOI22_X1 U12571 ( .A1(n16750), .A2(n12281), .B1(n16744), .B2(n16463), .ZN(
        n14071) );
  AOI22_X1 U12572 ( .A1(n16750), .A2(n12280), .B1(n16744), .B2(n16464), .ZN(
        n14053) );
  AOI22_X1 U12573 ( .A1(n16750), .A2(n12279), .B1(n16744), .B2(n16465), .ZN(
        n14035) );
  AOI22_X1 U12574 ( .A1(n16750), .A2(n12278), .B1(n16744), .B2(n16466), .ZN(
        n14017) );
  AOI22_X1 U12575 ( .A1(n16727), .A2(n12213), .B1(n16721), .B2(n12405), .ZN(
        n14000) );
  AOI22_X1 U12576 ( .A1(n16727), .A2(n12212), .B1(n16721), .B2(n12404), .ZN(
        n13982) );
  AOI22_X1 U12577 ( .A1(n16727), .A2(n12211), .B1(n16721), .B2(n12403), .ZN(
        n13964) );
  AOI22_X1 U12578 ( .A1(n16727), .A2(n12210), .B1(n16721), .B2(n12402), .ZN(
        n13946) );
  AOI22_X1 U12579 ( .A1(n16727), .A2(n12209), .B1(n16721), .B2(n12401), .ZN(
        n13928) );
  AOI22_X1 U12580 ( .A1(n16727), .A2(n12208), .B1(n16721), .B2(n12400), .ZN(
        n13910) );
  AOI22_X1 U12581 ( .A1(n16727), .A2(n12207), .B1(n16721), .B2(n12399), .ZN(
        n13892) );
  AOI22_X1 U12582 ( .A1(n16727), .A2(n12206), .B1(n16721), .B2(n12398), .ZN(
        n13874) );
  AOI22_X1 U12583 ( .A1(n16727), .A2(n12205), .B1(n16721), .B2(n12397), .ZN(
        n13856) );
  AOI22_X1 U12584 ( .A1(n16727), .A2(n12204), .B1(n16721), .B2(n12396), .ZN(
        n13838) );
  AOI22_X1 U12585 ( .A1(n16727), .A2(n12203), .B1(n16721), .B2(n12395), .ZN(
        n13820) );
  AOI22_X1 U12586 ( .A1(n16727), .A2(n12202), .B1(n16721), .B2(n12394), .ZN(
        n13802) );
  AOI22_X1 U12587 ( .A1(n16728), .A2(n12201), .B1(n16722), .B2(n12393), .ZN(
        n13784) );
  AOI22_X1 U12588 ( .A1(n16728), .A2(n12200), .B1(n16722), .B2(n12392), .ZN(
        n13766) );
  AOI22_X1 U12589 ( .A1(n16728), .A2(n12199), .B1(n16722), .B2(n12391), .ZN(
        n13748) );
  AOI22_X1 U12590 ( .A1(n16728), .A2(n12198), .B1(n16722), .B2(n12390), .ZN(
        n13723) );
  OAI22_X1 U12591 ( .A1(n16897), .A2(n17480), .B1(n16891), .B2(n13546), .ZN(
        n5028) );
  OAI22_X1 U12592 ( .A1(n16898), .A2(n17482), .B1(n16892), .B2(n13545), .ZN(
        n5029) );
  OAI22_X1 U12593 ( .A1(n16898), .A2(n17484), .B1(n16890), .B2(n13544), .ZN(
        n5030) );
  OAI22_X1 U12594 ( .A1(n16898), .A2(n17486), .B1(n16891), .B2(n13543), .ZN(
        n5031) );
  OAI22_X1 U12595 ( .A1(n16898), .A2(n17488), .B1(n16892), .B2(n13542), .ZN(
        n5032) );
  OAI22_X1 U12596 ( .A1(n16898), .A2(n17490), .B1(n16890), .B2(n13541), .ZN(
        n5033) );
  OAI22_X1 U12597 ( .A1(n16899), .A2(n17492), .B1(n16891), .B2(n13540), .ZN(
        n5034) );
  OAI22_X1 U12598 ( .A1(n16899), .A2(n17494), .B1(n16892), .B2(n13539), .ZN(
        n5035) );
  OAI22_X1 U12599 ( .A1(n16899), .A2(n17496), .B1(n16890), .B2(n13538), .ZN(
        n5036) );
  OAI22_X1 U12600 ( .A1(n16899), .A2(n17498), .B1(n16891), .B2(n13537), .ZN(
        n5037) );
  OAI22_X1 U12601 ( .A1(n16899), .A2(n17500), .B1(n16892), .B2(n13536), .ZN(
        n5038) );
  OAI22_X1 U12602 ( .A1(n16900), .A2(n17502), .B1(n16890), .B2(n13535), .ZN(
        n5039) );
  OAI22_X1 U12603 ( .A1(n16900), .A2(n17504), .B1(n13679), .B2(n13534), .ZN(
        n5040) );
  OAI22_X1 U12604 ( .A1(n16900), .A2(n17506), .B1(n16890), .B2(n13533), .ZN(
        n5041) );
  OAI22_X1 U12605 ( .A1(n16900), .A2(n17508), .B1(n13679), .B2(n13532), .ZN(
        n5042) );
  OAI22_X1 U12606 ( .A1(n16900), .A2(n17510), .B1(n16890), .B2(n13531), .ZN(
        n5043) );
  OAI22_X1 U12607 ( .A1(n16901), .A2(n17512), .B1(n13679), .B2(n13530), .ZN(
        n5044) );
  OAI22_X1 U12608 ( .A1(n16901), .A2(n17514), .B1(n16890), .B2(n13529), .ZN(
        n5045) );
  OAI22_X1 U12609 ( .A1(n16901), .A2(n17516), .B1(n16891), .B2(n13528), .ZN(
        n5046) );
  OAI22_X1 U12610 ( .A1(n16901), .A2(n17518), .B1(n16892), .B2(n13527), .ZN(
        n5047) );
  OAI22_X1 U12611 ( .A1(n16901), .A2(n17520), .B1(n16890), .B2(n13526), .ZN(
        n5048) );
  OAI22_X1 U12612 ( .A1(n16902), .A2(n17522), .B1(n16890), .B2(n13525), .ZN(
        n5049) );
  OAI22_X1 U12613 ( .A1(n16902), .A2(n17524), .B1(n16891), .B2(n13524), .ZN(
        n5050) );
  OAI22_X1 U12614 ( .A1(n16902), .A2(n17526), .B1(n16892), .B2(n13523), .ZN(
        n5051) );
  OAI22_X1 U12615 ( .A1(n16902), .A2(n17528), .B1(n16890), .B2(n13522), .ZN(
        n5052) );
  OAI22_X1 U12616 ( .A1(n16902), .A2(n17530), .B1(n16890), .B2(n13521), .ZN(
        n5053) );
  OAI22_X1 U12617 ( .A1(n16903), .A2(n17532), .B1(n13679), .B2(n13520), .ZN(
        n5054) );
  OAI22_X1 U12618 ( .A1(n16903), .A2(n17534), .B1(n16890), .B2(n13519), .ZN(
        n5055) );
  OAI22_X1 U12619 ( .A1(n16903), .A2(n17536), .B1(n13679), .B2(n13518), .ZN(
        n5056) );
  OAI22_X1 U12620 ( .A1(n16903), .A2(n17538), .B1(n16890), .B2(n13517), .ZN(
        n5057) );
  OAI22_X1 U12621 ( .A1(n16903), .A2(n17540), .B1(n13679), .B2(n13516), .ZN(
        n5058) );
  OAI22_X1 U12622 ( .A1(n16904), .A2(n17542), .B1(n16890), .B2(n13515), .ZN(
        n5059) );
  OAI22_X1 U12623 ( .A1(n16904), .A2(n17544), .B1(n13679), .B2(n13514), .ZN(
        n5060) );
  OAI22_X1 U12624 ( .A1(n16904), .A2(n17546), .B1(n16890), .B2(n13513), .ZN(
        n5061) );
  OAI22_X1 U12625 ( .A1(n16904), .A2(n17548), .B1(n13679), .B2(n13512), .ZN(
        n5062) );
  OAI22_X1 U12626 ( .A1(n16904), .A2(n17550), .B1(n16890), .B2(n13511), .ZN(
        n5063) );
  OAI22_X1 U12627 ( .A1(n16914), .A2(n17480), .B1(n16908), .B2(n13482), .ZN(
        n5092) );
  OAI22_X1 U12628 ( .A1(n16915), .A2(n17482), .B1(n16909), .B2(n13481), .ZN(
        n5093) );
  OAI22_X1 U12629 ( .A1(n16915), .A2(n17484), .B1(n16907), .B2(n13480), .ZN(
        n5094) );
  OAI22_X1 U12630 ( .A1(n16915), .A2(n17486), .B1(n16908), .B2(n13479), .ZN(
        n5095) );
  OAI22_X1 U12631 ( .A1(n16915), .A2(n17488), .B1(n16909), .B2(n13478), .ZN(
        n5096) );
  OAI22_X1 U12632 ( .A1(n16915), .A2(n17490), .B1(n16907), .B2(n13477), .ZN(
        n5097) );
  OAI22_X1 U12633 ( .A1(n16916), .A2(n17492), .B1(n16908), .B2(n13476), .ZN(
        n5098) );
  OAI22_X1 U12634 ( .A1(n16916), .A2(n17494), .B1(n16909), .B2(n13475), .ZN(
        n5099) );
  OAI22_X1 U12635 ( .A1(n16916), .A2(n17496), .B1(n16907), .B2(n13474), .ZN(
        n5100) );
  OAI22_X1 U12636 ( .A1(n16916), .A2(n17498), .B1(n16908), .B2(n13473), .ZN(
        n5101) );
  OAI22_X1 U12637 ( .A1(n16916), .A2(n17500), .B1(n16909), .B2(n13472), .ZN(
        n5102) );
  OAI22_X1 U12638 ( .A1(n16917), .A2(n17502), .B1(n16907), .B2(n13471), .ZN(
        n5103) );
  OAI22_X1 U12639 ( .A1(n16917), .A2(n17504), .B1(n13678), .B2(n13470), .ZN(
        n5104) );
  OAI22_X1 U12640 ( .A1(n16917), .A2(n17506), .B1(n16907), .B2(n13469), .ZN(
        n5105) );
  OAI22_X1 U12641 ( .A1(n16917), .A2(n17508), .B1(n13678), .B2(n13468), .ZN(
        n5106) );
  OAI22_X1 U12642 ( .A1(n16917), .A2(n17510), .B1(n16907), .B2(n13467), .ZN(
        n5107) );
  OAI22_X1 U12643 ( .A1(n16918), .A2(n17512), .B1(n13678), .B2(n13466), .ZN(
        n5108) );
  OAI22_X1 U12644 ( .A1(n16918), .A2(n17514), .B1(n16907), .B2(n13465), .ZN(
        n5109) );
  OAI22_X1 U12645 ( .A1(n16918), .A2(n17516), .B1(n16908), .B2(n13464), .ZN(
        n5110) );
  OAI22_X1 U12646 ( .A1(n16918), .A2(n17518), .B1(n16909), .B2(n13463), .ZN(
        n5111) );
  OAI22_X1 U12647 ( .A1(n16918), .A2(n17520), .B1(n16907), .B2(n13462), .ZN(
        n5112) );
  OAI22_X1 U12648 ( .A1(n16919), .A2(n17522), .B1(n16907), .B2(n13461), .ZN(
        n5113) );
  OAI22_X1 U12649 ( .A1(n16919), .A2(n17524), .B1(n16908), .B2(n13460), .ZN(
        n5114) );
  OAI22_X1 U12650 ( .A1(n16919), .A2(n17526), .B1(n16909), .B2(n13459), .ZN(
        n5115) );
  OAI22_X1 U12651 ( .A1(n16919), .A2(n17528), .B1(n16907), .B2(n13458), .ZN(
        n5116) );
  OAI22_X1 U12652 ( .A1(n16919), .A2(n17530), .B1(n16907), .B2(n13457), .ZN(
        n5117) );
  OAI22_X1 U12653 ( .A1(n16920), .A2(n17532), .B1(n13678), .B2(n13456), .ZN(
        n5118) );
  OAI22_X1 U12654 ( .A1(n16920), .A2(n17534), .B1(n16907), .B2(n13455), .ZN(
        n5119) );
  OAI22_X1 U12655 ( .A1(n16920), .A2(n17536), .B1(n13678), .B2(n13454), .ZN(
        n5120) );
  OAI22_X1 U12656 ( .A1(n16920), .A2(n17538), .B1(n16907), .B2(n13453), .ZN(
        n5121) );
  OAI22_X1 U12657 ( .A1(n16920), .A2(n17540), .B1(n13678), .B2(n13452), .ZN(
        n5122) );
  OAI22_X1 U12658 ( .A1(n16921), .A2(n17542), .B1(n16907), .B2(n13451), .ZN(
        n5123) );
  OAI22_X1 U12659 ( .A1(n16921), .A2(n17544), .B1(n13678), .B2(n13450), .ZN(
        n5124) );
  OAI22_X1 U12660 ( .A1(n16921), .A2(n17546), .B1(n16907), .B2(n13449), .ZN(
        n5125) );
  OAI22_X1 U12661 ( .A1(n16921), .A2(n17548), .B1(n13678), .B2(n13448), .ZN(
        n5126) );
  OAI22_X1 U12662 ( .A1(n16921), .A2(n17550), .B1(n16907), .B2(n13447), .ZN(
        n5127) );
  OAI22_X1 U12663 ( .A1(n17067), .A2(n17480), .B1(n17061), .B2(n13034), .ZN(
        n5668) );
  OAI22_X1 U12664 ( .A1(n17068), .A2(n17482), .B1(n17062), .B2(n13033), .ZN(
        n5669) );
  OAI22_X1 U12665 ( .A1(n17068), .A2(n17484), .B1(n17060), .B2(n13032), .ZN(
        n5670) );
  OAI22_X1 U12666 ( .A1(n17068), .A2(n17486), .B1(n17061), .B2(n13031), .ZN(
        n5671) );
  OAI22_X1 U12667 ( .A1(n17068), .A2(n17488), .B1(n17062), .B2(n13030), .ZN(
        n5672) );
  OAI22_X1 U12668 ( .A1(n17068), .A2(n17490), .B1(n17060), .B2(n13029), .ZN(
        n5673) );
  OAI22_X1 U12669 ( .A1(n17069), .A2(n17492), .B1(n17061), .B2(n13028), .ZN(
        n5674) );
  OAI22_X1 U12670 ( .A1(n17069), .A2(n17494), .B1(n17062), .B2(n13027), .ZN(
        n5675) );
  OAI22_X1 U12671 ( .A1(n17069), .A2(n17496), .B1(n17060), .B2(n13026), .ZN(
        n5676) );
  OAI22_X1 U12672 ( .A1(n17069), .A2(n17498), .B1(n17061), .B2(n13025), .ZN(
        n5677) );
  OAI22_X1 U12673 ( .A1(n17069), .A2(n17500), .B1(n17062), .B2(n13024), .ZN(
        n5678) );
  OAI22_X1 U12674 ( .A1(n17070), .A2(n17502), .B1(n17060), .B2(n13023), .ZN(
        n5679) );
  OAI22_X1 U12675 ( .A1(n17070), .A2(n17504), .B1(n13668), .B2(n13022), .ZN(
        n5680) );
  OAI22_X1 U12676 ( .A1(n17070), .A2(n17506), .B1(n17060), .B2(n13021), .ZN(
        n5681) );
  OAI22_X1 U12677 ( .A1(n17070), .A2(n17508), .B1(n13668), .B2(n13020), .ZN(
        n5682) );
  OAI22_X1 U12678 ( .A1(n17070), .A2(n17510), .B1(n17060), .B2(n13019), .ZN(
        n5683) );
  OAI22_X1 U12679 ( .A1(n17071), .A2(n17512), .B1(n13668), .B2(n13018), .ZN(
        n5684) );
  OAI22_X1 U12680 ( .A1(n17071), .A2(n17514), .B1(n17060), .B2(n13017), .ZN(
        n5685) );
  OAI22_X1 U12681 ( .A1(n17071), .A2(n17516), .B1(n17061), .B2(n13016), .ZN(
        n5686) );
  OAI22_X1 U12682 ( .A1(n17071), .A2(n17518), .B1(n17062), .B2(n13015), .ZN(
        n5687) );
  OAI22_X1 U12683 ( .A1(n17071), .A2(n17520), .B1(n17060), .B2(n13014), .ZN(
        n5688) );
  OAI22_X1 U12684 ( .A1(n17072), .A2(n17522), .B1(n17060), .B2(n13013), .ZN(
        n5689) );
  OAI22_X1 U12685 ( .A1(n17072), .A2(n17524), .B1(n17061), .B2(n13012), .ZN(
        n5690) );
  OAI22_X1 U12686 ( .A1(n17072), .A2(n17526), .B1(n17062), .B2(n13011), .ZN(
        n5691) );
  OAI22_X1 U12687 ( .A1(n17072), .A2(n17528), .B1(n17060), .B2(n13010), .ZN(
        n5692) );
  OAI22_X1 U12688 ( .A1(n17072), .A2(n17530), .B1(n17060), .B2(n13009), .ZN(
        n5693) );
  OAI22_X1 U12689 ( .A1(n17073), .A2(n17532), .B1(n13668), .B2(n13008), .ZN(
        n5694) );
  OAI22_X1 U12690 ( .A1(n17073), .A2(n17534), .B1(n17060), .B2(n13007), .ZN(
        n5695) );
  OAI22_X1 U12691 ( .A1(n17073), .A2(n17536), .B1(n13668), .B2(n13006), .ZN(
        n5696) );
  OAI22_X1 U12692 ( .A1(n17073), .A2(n17538), .B1(n17060), .B2(n13005), .ZN(
        n5697) );
  OAI22_X1 U12693 ( .A1(n17073), .A2(n17540), .B1(n13668), .B2(n13004), .ZN(
        n5698) );
  OAI22_X1 U12694 ( .A1(n17074), .A2(n17542), .B1(n17060), .B2(n13003), .ZN(
        n5699) );
  OAI22_X1 U12695 ( .A1(n17074), .A2(n17544), .B1(n13668), .B2(n13002), .ZN(
        n5700) );
  OAI22_X1 U12696 ( .A1(n17074), .A2(n17546), .B1(n17060), .B2(n13001), .ZN(
        n5701) );
  OAI22_X1 U12697 ( .A1(n17074), .A2(n17548), .B1(n13668), .B2(n13000), .ZN(
        n5702) );
  OAI22_X1 U12698 ( .A1(n17074), .A2(n17550), .B1(n17060), .B2(n12999), .ZN(
        n5703) );
  OAI22_X1 U12699 ( .A1(n17221), .A2(n17481), .B1(n17215), .B2(n12749), .ZN(
        n6244) );
  OAI22_X1 U12700 ( .A1(n17222), .A2(n17483), .B1(n17216), .B2(n12748), .ZN(
        n6245) );
  OAI22_X1 U12701 ( .A1(n17222), .A2(n17485), .B1(n17214), .B2(n12747), .ZN(
        n6246) );
  OAI22_X1 U12702 ( .A1(n17222), .A2(n17487), .B1(n17215), .B2(n12746), .ZN(
        n6247) );
  OAI22_X1 U12703 ( .A1(n17222), .A2(n17489), .B1(n17216), .B2(n12745), .ZN(
        n6248) );
  OAI22_X1 U12704 ( .A1(n17222), .A2(n17491), .B1(n17214), .B2(n12744), .ZN(
        n6249) );
  OAI22_X1 U12705 ( .A1(n17223), .A2(n17493), .B1(n17215), .B2(n12743), .ZN(
        n6250) );
  OAI22_X1 U12706 ( .A1(n17223), .A2(n17495), .B1(n17216), .B2(n12742), .ZN(
        n6251) );
  OAI22_X1 U12707 ( .A1(n17223), .A2(n17497), .B1(n17214), .B2(n12741), .ZN(
        n6252) );
  OAI22_X1 U12708 ( .A1(n17223), .A2(n17499), .B1(n17215), .B2(n12740), .ZN(
        n6253) );
  OAI22_X1 U12709 ( .A1(n17223), .A2(n17501), .B1(n17216), .B2(n12739), .ZN(
        n6254) );
  OAI22_X1 U12710 ( .A1(n17224), .A2(n17503), .B1(n17214), .B2(n12738), .ZN(
        n6255) );
  OAI22_X1 U12711 ( .A1(n17224), .A2(n17505), .B1(n13658), .B2(n12737), .ZN(
        n6256) );
  OAI22_X1 U12712 ( .A1(n17224), .A2(n17507), .B1(n17214), .B2(n12736), .ZN(
        n6257) );
  OAI22_X1 U12713 ( .A1(n17224), .A2(n17509), .B1(n13658), .B2(n12735), .ZN(
        n6258) );
  OAI22_X1 U12714 ( .A1(n17224), .A2(n17511), .B1(n17214), .B2(n12734), .ZN(
        n6259) );
  OAI22_X1 U12715 ( .A1(n17225), .A2(n17513), .B1(n13658), .B2(n12733), .ZN(
        n6260) );
  OAI22_X1 U12716 ( .A1(n17225), .A2(n17515), .B1(n17214), .B2(n12732), .ZN(
        n6261) );
  OAI22_X1 U12717 ( .A1(n17225), .A2(n17517), .B1(n17215), .B2(n12731), .ZN(
        n6262) );
  OAI22_X1 U12718 ( .A1(n17225), .A2(n17519), .B1(n17216), .B2(n12730), .ZN(
        n6263) );
  OAI22_X1 U12719 ( .A1(n17225), .A2(n17521), .B1(n17214), .B2(n12729), .ZN(
        n6264) );
  OAI22_X1 U12720 ( .A1(n17226), .A2(n17523), .B1(n17214), .B2(n12728), .ZN(
        n6265) );
  OAI22_X1 U12721 ( .A1(n17226), .A2(n17525), .B1(n17215), .B2(n12727), .ZN(
        n6266) );
  OAI22_X1 U12722 ( .A1(n17226), .A2(n17527), .B1(n17216), .B2(n12726), .ZN(
        n6267) );
  OAI22_X1 U12723 ( .A1(n17226), .A2(n17529), .B1(n17214), .B2(n12725), .ZN(
        n6268) );
  OAI22_X1 U12724 ( .A1(n17226), .A2(n17531), .B1(n17214), .B2(n12724), .ZN(
        n6269) );
  OAI22_X1 U12725 ( .A1(n17227), .A2(n17533), .B1(n13658), .B2(n12723), .ZN(
        n6270) );
  OAI22_X1 U12726 ( .A1(n17227), .A2(n17535), .B1(n17214), .B2(n12722), .ZN(
        n6271) );
  OAI22_X1 U12727 ( .A1(n17227), .A2(n17537), .B1(n13658), .B2(n12721), .ZN(
        n6272) );
  OAI22_X1 U12728 ( .A1(n17227), .A2(n17539), .B1(n17214), .B2(n12720), .ZN(
        n6273) );
  OAI22_X1 U12729 ( .A1(n17227), .A2(n17541), .B1(n13658), .B2(n12719), .ZN(
        n6274) );
  OAI22_X1 U12730 ( .A1(n17228), .A2(n17543), .B1(n17214), .B2(n12718), .ZN(
        n6275) );
  OAI22_X1 U12731 ( .A1(n17228), .A2(n17545), .B1(n13658), .B2(n12717), .ZN(
        n6276) );
  OAI22_X1 U12732 ( .A1(n17228), .A2(n17547), .B1(n17214), .B2(n12716), .ZN(
        n6277) );
  OAI22_X1 U12733 ( .A1(n17228), .A2(n17549), .B1(n13658), .B2(n12715), .ZN(
        n6278) );
  OAI22_X1 U12734 ( .A1(n17228), .A2(n17551), .B1(n17214), .B2(n12714), .ZN(
        n6279) );
  OAI22_X1 U12735 ( .A1(n17255), .A2(n17481), .B1(n17249), .B2(n12621), .ZN(
        n6372) );
  OAI22_X1 U12736 ( .A1(n17256), .A2(n17483), .B1(n17250), .B2(n12620), .ZN(
        n6373) );
  OAI22_X1 U12737 ( .A1(n17256), .A2(n17485), .B1(n17248), .B2(n12619), .ZN(
        n6374) );
  OAI22_X1 U12738 ( .A1(n17256), .A2(n17487), .B1(n17249), .B2(n12618), .ZN(
        n6375) );
  OAI22_X1 U12739 ( .A1(n17256), .A2(n17489), .B1(n17250), .B2(n12617), .ZN(
        n6376) );
  OAI22_X1 U12740 ( .A1(n17256), .A2(n17491), .B1(n17248), .B2(n12616), .ZN(
        n6377) );
  OAI22_X1 U12741 ( .A1(n17257), .A2(n17493), .B1(n17249), .B2(n12615), .ZN(
        n6378) );
  OAI22_X1 U12742 ( .A1(n17257), .A2(n17495), .B1(n17250), .B2(n12614), .ZN(
        n6379) );
  OAI22_X1 U12743 ( .A1(n17257), .A2(n17497), .B1(n17248), .B2(n12613), .ZN(
        n6380) );
  OAI22_X1 U12744 ( .A1(n17257), .A2(n17499), .B1(n17249), .B2(n12612), .ZN(
        n6381) );
  OAI22_X1 U12745 ( .A1(n17257), .A2(n17501), .B1(n17250), .B2(n12611), .ZN(
        n6382) );
  OAI22_X1 U12746 ( .A1(n17258), .A2(n17503), .B1(n17248), .B2(n12610), .ZN(
        n6383) );
  OAI22_X1 U12747 ( .A1(n17258), .A2(n17505), .B1(n13656), .B2(n12609), .ZN(
        n6384) );
  OAI22_X1 U12748 ( .A1(n17258), .A2(n17507), .B1(n17248), .B2(n12608), .ZN(
        n6385) );
  OAI22_X1 U12749 ( .A1(n17258), .A2(n17509), .B1(n13656), .B2(n12607), .ZN(
        n6386) );
  OAI22_X1 U12750 ( .A1(n17258), .A2(n17511), .B1(n17248), .B2(n12606), .ZN(
        n6387) );
  OAI22_X1 U12751 ( .A1(n17259), .A2(n17513), .B1(n13656), .B2(n12605), .ZN(
        n6388) );
  OAI22_X1 U12752 ( .A1(n17259), .A2(n17515), .B1(n17248), .B2(n12604), .ZN(
        n6389) );
  OAI22_X1 U12753 ( .A1(n17259), .A2(n17517), .B1(n17249), .B2(n12603), .ZN(
        n6390) );
  OAI22_X1 U12754 ( .A1(n17259), .A2(n17519), .B1(n17250), .B2(n12602), .ZN(
        n6391) );
  OAI22_X1 U12755 ( .A1(n17259), .A2(n17521), .B1(n17248), .B2(n12601), .ZN(
        n6392) );
  OAI22_X1 U12756 ( .A1(n17260), .A2(n17523), .B1(n17248), .B2(n12600), .ZN(
        n6393) );
  OAI22_X1 U12757 ( .A1(n17260), .A2(n17525), .B1(n17249), .B2(n12599), .ZN(
        n6394) );
  OAI22_X1 U12758 ( .A1(n17260), .A2(n17527), .B1(n17250), .B2(n12598), .ZN(
        n6395) );
  OAI22_X1 U12759 ( .A1(n17260), .A2(n17529), .B1(n17248), .B2(n12597), .ZN(
        n6396) );
  OAI22_X1 U12760 ( .A1(n17260), .A2(n17531), .B1(n17248), .B2(n12596), .ZN(
        n6397) );
  OAI22_X1 U12761 ( .A1(n17261), .A2(n17533), .B1(n13656), .B2(n12595), .ZN(
        n6398) );
  OAI22_X1 U12762 ( .A1(n17261), .A2(n17535), .B1(n17248), .B2(n12594), .ZN(
        n6399) );
  OAI22_X1 U12763 ( .A1(n17261), .A2(n17537), .B1(n13656), .B2(n12593), .ZN(
        n6400) );
  OAI22_X1 U12764 ( .A1(n17261), .A2(n17539), .B1(n17248), .B2(n12592), .ZN(
        n6401) );
  OAI22_X1 U12765 ( .A1(n17261), .A2(n17541), .B1(n13656), .B2(n12591), .ZN(
        n6402) );
  OAI22_X1 U12766 ( .A1(n17262), .A2(n17543), .B1(n17248), .B2(n12590), .ZN(
        n6403) );
  OAI22_X1 U12767 ( .A1(n17262), .A2(n17545), .B1(n13656), .B2(n12589), .ZN(
        n6404) );
  OAI22_X1 U12768 ( .A1(n17262), .A2(n17547), .B1(n17248), .B2(n12588), .ZN(
        n6405) );
  OAI22_X1 U12769 ( .A1(n17262), .A2(n17549), .B1(n13656), .B2(n12587), .ZN(
        n6406) );
  OAI22_X1 U12770 ( .A1(n17262), .A2(n17551), .B1(n17248), .B2(n12586), .ZN(
        n6407) );
  OAI22_X1 U12771 ( .A1(n16905), .A2(n17552), .B1(n13679), .B2(n13510), .ZN(
        n5064) );
  OAI22_X1 U12772 ( .A1(n16905), .A2(n17554), .B1(n13679), .B2(n13509), .ZN(
        n5065) );
  OAI22_X1 U12773 ( .A1(n16905), .A2(n17556), .B1(n16890), .B2(n13508), .ZN(
        n5066) );
  OAI22_X1 U12774 ( .A1(n16905), .A2(n17577), .B1(n13679), .B2(n13507), .ZN(
        n5067) );
  OAI22_X1 U12775 ( .A1(n16922), .A2(n17552), .B1(n13678), .B2(n13446), .ZN(
        n5128) );
  OAI22_X1 U12776 ( .A1(n16922), .A2(n17554), .B1(n13678), .B2(n13445), .ZN(
        n5129) );
  OAI22_X1 U12777 ( .A1(n16922), .A2(n17556), .B1(n16907), .B2(n13444), .ZN(
        n5130) );
  OAI22_X1 U12778 ( .A1(n16922), .A2(n17577), .B1(n13678), .B2(n13443), .ZN(
        n5131) );
  OAI22_X1 U12779 ( .A1(n17075), .A2(n17552), .B1(n13668), .B2(n12998), .ZN(
        n5704) );
  OAI22_X1 U12780 ( .A1(n17075), .A2(n17554), .B1(n13668), .B2(n12997), .ZN(
        n5705) );
  OAI22_X1 U12781 ( .A1(n17075), .A2(n17556), .B1(n17060), .B2(n12996), .ZN(
        n5706) );
  OAI22_X1 U12782 ( .A1(n17075), .A2(n17577), .B1(n13668), .B2(n12995), .ZN(
        n5707) );
  OAI22_X1 U12783 ( .A1(n17165), .A2(n17433), .B1(n13661), .B2(n12802), .ZN(
        n6028) );
  OAI22_X1 U12784 ( .A1(n17165), .A2(n17435), .B1(n13661), .B2(n12801), .ZN(
        n6029) );
  OAI22_X1 U12785 ( .A1(n17229), .A2(n17553), .B1(n13658), .B2(n12713), .ZN(
        n6280) );
  OAI22_X1 U12786 ( .A1(n17229), .A2(n17555), .B1(n13658), .B2(n12712), .ZN(
        n6281) );
  OAI22_X1 U12787 ( .A1(n17229), .A2(n17557), .B1(n17214), .B2(n12711), .ZN(
        n6282) );
  OAI22_X1 U12788 ( .A1(n17229), .A2(n17578), .B1(n13658), .B2(n12710), .ZN(
        n6283) );
  OAI22_X1 U12789 ( .A1(n17263), .A2(n17553), .B1(n13656), .B2(n12585), .ZN(
        n6408) );
  OAI22_X1 U12790 ( .A1(n17263), .A2(n17555), .B1(n13656), .B2(n12584), .ZN(
        n6409) );
  OAI22_X1 U12791 ( .A1(n17263), .A2(n17557), .B1(n17248), .B2(n12583), .ZN(
        n6410) );
  OAI22_X1 U12792 ( .A1(n17263), .A2(n17578), .B1(n13656), .B2(n12582), .ZN(
        n6411) );
  NAND2_X1 U12793 ( .A1(n16038), .A2(n16039), .ZN(n4877) );
  NOR4_X1 U12794 ( .A1(n16048), .A2(n16049), .A3(n16050), .A4(n16051), .ZN(
        n16038) );
  NOR4_X1 U12795 ( .A1(n16040), .A2(n16041), .A3(n16042), .A4(n16043), .ZN(
        n16039) );
  OAI221_X1 U12796 ( .B1(n13505), .B2(n16530), .C1(n12801), .C2(n16524), .A(
        n16054), .ZN(n16049) );
  NAND2_X1 U12797 ( .A1(n16020), .A2(n16021), .ZN(n4878) );
  NOR4_X1 U12798 ( .A1(n16030), .A2(n16031), .A3(n16032), .A4(n16033), .ZN(
        n16020) );
  NOR4_X1 U12799 ( .A1(n16022), .A2(n16023), .A3(n16024), .A4(n16025), .ZN(
        n16021) );
  OAI221_X1 U12800 ( .B1(n13504), .B2(n16530), .C1(n12800), .C2(n16524), .A(
        n16036), .ZN(n16031) );
  NAND2_X1 U12801 ( .A1(n16002), .A2(n16003), .ZN(n4879) );
  NOR4_X1 U12802 ( .A1(n16012), .A2(n16013), .A3(n16014), .A4(n16015), .ZN(
        n16002) );
  NOR4_X1 U12803 ( .A1(n16004), .A2(n16005), .A3(n16006), .A4(n16007), .ZN(
        n16003) );
  OAI221_X1 U12804 ( .B1(n13503), .B2(n16530), .C1(n12799), .C2(n16524), .A(
        n16018), .ZN(n16013) );
  NAND2_X1 U12805 ( .A1(n15984), .A2(n15985), .ZN(n4880) );
  NOR4_X1 U12806 ( .A1(n15994), .A2(n15995), .A3(n15996), .A4(n15997), .ZN(
        n15984) );
  NOR4_X1 U12807 ( .A1(n15986), .A2(n15987), .A3(n15988), .A4(n15989), .ZN(
        n15985) );
  OAI221_X1 U12808 ( .B1(n13502), .B2(n16530), .C1(n12798), .C2(n16524), .A(
        n16000), .ZN(n15995) );
  NAND2_X1 U12809 ( .A1(n15966), .A2(n15967), .ZN(n4881) );
  NOR4_X1 U12810 ( .A1(n15976), .A2(n15977), .A3(n15978), .A4(n15979), .ZN(
        n15966) );
  NOR4_X1 U12811 ( .A1(n15968), .A2(n15969), .A3(n15970), .A4(n15971), .ZN(
        n15967) );
  OAI221_X1 U12812 ( .B1(n13501), .B2(n16530), .C1(n12797), .C2(n16524), .A(
        n15982), .ZN(n15977) );
  NAND2_X1 U12813 ( .A1(n15948), .A2(n15949), .ZN(n4882) );
  NOR4_X1 U12814 ( .A1(n15958), .A2(n15959), .A3(n15960), .A4(n15961), .ZN(
        n15948) );
  NOR4_X1 U12815 ( .A1(n15950), .A2(n15951), .A3(n15952), .A4(n15953), .ZN(
        n15949) );
  OAI221_X1 U12816 ( .B1(n13500), .B2(n16530), .C1(n12796), .C2(n16524), .A(
        n15964), .ZN(n15959) );
  NAND2_X1 U12817 ( .A1(n15930), .A2(n15931), .ZN(n4883) );
  NOR4_X1 U12818 ( .A1(n15940), .A2(n15941), .A3(n15942), .A4(n15943), .ZN(
        n15930) );
  NOR4_X1 U12819 ( .A1(n15932), .A2(n15933), .A3(n15934), .A4(n15935), .ZN(
        n15931) );
  OAI221_X1 U12820 ( .B1(n13499), .B2(n16530), .C1(n12795), .C2(n16524), .A(
        n15946), .ZN(n15941) );
  NAND2_X1 U12821 ( .A1(n15912), .A2(n15913), .ZN(n4884) );
  NOR4_X1 U12822 ( .A1(n15922), .A2(n15923), .A3(n15924), .A4(n15925), .ZN(
        n15912) );
  NOR4_X1 U12823 ( .A1(n15914), .A2(n15915), .A3(n15916), .A4(n15917), .ZN(
        n15913) );
  OAI221_X1 U12824 ( .B1(n13498), .B2(n16530), .C1(n12794), .C2(n16524), .A(
        n15928), .ZN(n15923) );
  NAND2_X1 U12825 ( .A1(n15894), .A2(n15895), .ZN(n4885) );
  NOR4_X1 U12826 ( .A1(n15904), .A2(n15905), .A3(n15906), .A4(n15907), .ZN(
        n15894) );
  NOR4_X1 U12827 ( .A1(n15896), .A2(n15897), .A3(n15898), .A4(n15899), .ZN(
        n15895) );
  OAI221_X1 U12828 ( .B1(n13497), .B2(n16530), .C1(n12793), .C2(n16524), .A(
        n15910), .ZN(n15905) );
  NAND2_X1 U12829 ( .A1(n15876), .A2(n15877), .ZN(n4886) );
  NOR4_X1 U12830 ( .A1(n15886), .A2(n15887), .A3(n15888), .A4(n15889), .ZN(
        n15876) );
  NOR4_X1 U12831 ( .A1(n15878), .A2(n15879), .A3(n15880), .A4(n15881), .ZN(
        n15877) );
  OAI221_X1 U12832 ( .B1(n13496), .B2(n16530), .C1(n12792), .C2(n16524), .A(
        n15892), .ZN(n15887) );
  NAND2_X1 U12833 ( .A1(n15858), .A2(n15859), .ZN(n4887) );
  NOR4_X1 U12834 ( .A1(n15868), .A2(n15869), .A3(n15870), .A4(n15871), .ZN(
        n15858) );
  NOR4_X1 U12835 ( .A1(n15860), .A2(n15861), .A3(n15862), .A4(n15863), .ZN(
        n15859) );
  OAI221_X1 U12836 ( .B1(n13495), .B2(n16530), .C1(n12791), .C2(n16524), .A(
        n15874), .ZN(n15869) );
  NAND2_X1 U12837 ( .A1(n15840), .A2(n15841), .ZN(n4888) );
  NOR4_X1 U12838 ( .A1(n15850), .A2(n15851), .A3(n15852), .A4(n15853), .ZN(
        n15840) );
  NOR4_X1 U12839 ( .A1(n15842), .A2(n15843), .A3(n15844), .A4(n15845), .ZN(
        n15841) );
  OAI221_X1 U12840 ( .B1(n13494), .B2(n16531), .C1(n12790), .C2(n16525), .A(
        n15856), .ZN(n15851) );
  NAND2_X1 U12841 ( .A1(n15822), .A2(n15823), .ZN(n4889) );
  NOR4_X1 U12842 ( .A1(n15832), .A2(n15833), .A3(n15834), .A4(n15835), .ZN(
        n15822) );
  NOR4_X1 U12843 ( .A1(n15824), .A2(n15825), .A3(n15826), .A4(n15827), .ZN(
        n15823) );
  OAI221_X1 U12844 ( .B1(n13493), .B2(n16531), .C1(n12789), .C2(n16525), .A(
        n15838), .ZN(n15833) );
  NAND2_X1 U12845 ( .A1(n15804), .A2(n15805), .ZN(n4890) );
  NOR4_X1 U12846 ( .A1(n15814), .A2(n15815), .A3(n15816), .A4(n15817), .ZN(
        n15804) );
  NOR4_X1 U12847 ( .A1(n15806), .A2(n15807), .A3(n15808), .A4(n15809), .ZN(
        n15805) );
  OAI221_X1 U12848 ( .B1(n13492), .B2(n16531), .C1(n12788), .C2(n16525), .A(
        n15820), .ZN(n15815) );
  NAND2_X1 U12849 ( .A1(n15786), .A2(n15787), .ZN(n4891) );
  NOR4_X1 U12850 ( .A1(n15796), .A2(n15797), .A3(n15798), .A4(n15799), .ZN(
        n15786) );
  NOR4_X1 U12851 ( .A1(n15788), .A2(n15789), .A3(n15790), .A4(n15791), .ZN(
        n15787) );
  OAI221_X1 U12852 ( .B1(n13491), .B2(n16531), .C1(n12787), .C2(n16525), .A(
        n15802), .ZN(n15797) );
  NAND2_X1 U12853 ( .A1(n15768), .A2(n15769), .ZN(n4892) );
  NOR4_X1 U12854 ( .A1(n15778), .A2(n15779), .A3(n15780), .A4(n15781), .ZN(
        n15768) );
  NOR4_X1 U12855 ( .A1(n15770), .A2(n15771), .A3(n15772), .A4(n15773), .ZN(
        n15769) );
  OAI221_X1 U12856 ( .B1(n13490), .B2(n16531), .C1(n12786), .C2(n16525), .A(
        n15784), .ZN(n15779) );
  NAND2_X1 U12857 ( .A1(n15750), .A2(n15751), .ZN(n4893) );
  NOR4_X1 U12858 ( .A1(n15760), .A2(n15761), .A3(n15762), .A4(n15763), .ZN(
        n15750) );
  NOR4_X1 U12859 ( .A1(n15752), .A2(n15753), .A3(n15754), .A4(n15755), .ZN(
        n15751) );
  OAI221_X1 U12860 ( .B1(n13489), .B2(n16531), .C1(n12785), .C2(n16525), .A(
        n15766), .ZN(n15761) );
  NAND2_X1 U12861 ( .A1(n15732), .A2(n15733), .ZN(n4894) );
  NOR4_X1 U12862 ( .A1(n15742), .A2(n15743), .A3(n15744), .A4(n15745), .ZN(
        n15732) );
  NOR4_X1 U12863 ( .A1(n15734), .A2(n15735), .A3(n15736), .A4(n15737), .ZN(
        n15733) );
  OAI221_X1 U12864 ( .B1(n13488), .B2(n16531), .C1(n12784), .C2(n16525), .A(
        n15748), .ZN(n15743) );
  NAND2_X1 U12865 ( .A1(n15714), .A2(n15715), .ZN(n4895) );
  NOR4_X1 U12866 ( .A1(n15724), .A2(n15725), .A3(n15726), .A4(n15727), .ZN(
        n15714) );
  NOR4_X1 U12867 ( .A1(n15716), .A2(n15717), .A3(n15718), .A4(n15719), .ZN(
        n15715) );
  OAI221_X1 U12868 ( .B1(n13487), .B2(n16531), .C1(n12783), .C2(n16525), .A(
        n15730), .ZN(n15725) );
  NAND2_X1 U12869 ( .A1(n15696), .A2(n15697), .ZN(n4896) );
  NOR4_X1 U12870 ( .A1(n15706), .A2(n15707), .A3(n15708), .A4(n15709), .ZN(
        n15696) );
  NOR4_X1 U12871 ( .A1(n15698), .A2(n15699), .A3(n15700), .A4(n15701), .ZN(
        n15697) );
  OAI221_X1 U12872 ( .B1(n13486), .B2(n16531), .C1(n12782), .C2(n16525), .A(
        n15712), .ZN(n15707) );
  NAND2_X1 U12873 ( .A1(n15678), .A2(n15679), .ZN(n4897) );
  NOR4_X1 U12874 ( .A1(n15688), .A2(n15689), .A3(n15690), .A4(n15691), .ZN(
        n15678) );
  NOR4_X1 U12875 ( .A1(n15680), .A2(n15681), .A3(n15682), .A4(n15683), .ZN(
        n15679) );
  OAI221_X1 U12876 ( .B1(n13485), .B2(n16531), .C1(n12781), .C2(n16525), .A(
        n15694), .ZN(n15689) );
  NAND2_X1 U12877 ( .A1(n15660), .A2(n15661), .ZN(n4898) );
  NOR4_X1 U12878 ( .A1(n15670), .A2(n15671), .A3(n15672), .A4(n15673), .ZN(
        n15660) );
  NOR4_X1 U12879 ( .A1(n15662), .A2(n15663), .A3(n15664), .A4(n15665), .ZN(
        n15661) );
  OAI221_X1 U12880 ( .B1(n13484), .B2(n16531), .C1(n12780), .C2(n16525), .A(
        n15676), .ZN(n15671) );
  NAND2_X1 U12881 ( .A1(n15642), .A2(n15643), .ZN(n4899) );
  NOR4_X1 U12882 ( .A1(n15652), .A2(n15653), .A3(n15654), .A4(n15655), .ZN(
        n15642) );
  NOR4_X1 U12883 ( .A1(n15644), .A2(n15645), .A3(n15646), .A4(n15647), .ZN(
        n15643) );
  OAI221_X1 U12884 ( .B1(n13483), .B2(n16531), .C1(n12779), .C2(n16525), .A(
        n15658), .ZN(n15653) );
  NAND2_X1 U12885 ( .A1(n15624), .A2(n15625), .ZN(n4900) );
  NOR4_X1 U12886 ( .A1(n15634), .A2(n15635), .A3(n15636), .A4(n15637), .ZN(
        n15624) );
  NOR4_X1 U12887 ( .A1(n15626), .A2(n15627), .A3(n15628), .A4(n15629), .ZN(
        n15625) );
  OAI221_X1 U12888 ( .B1(n13482), .B2(n16532), .C1(n12778), .C2(n16526), .A(
        n15640), .ZN(n15635) );
  NAND2_X1 U12889 ( .A1(n15606), .A2(n15607), .ZN(n4901) );
  NOR4_X1 U12890 ( .A1(n15616), .A2(n15617), .A3(n15618), .A4(n15619), .ZN(
        n15606) );
  NOR4_X1 U12891 ( .A1(n15608), .A2(n15609), .A3(n15610), .A4(n15611), .ZN(
        n15607) );
  OAI221_X1 U12892 ( .B1(n13481), .B2(n16532), .C1(n12777), .C2(n16526), .A(
        n15622), .ZN(n15617) );
  NAND2_X1 U12893 ( .A1(n15588), .A2(n15589), .ZN(n4902) );
  NOR4_X1 U12894 ( .A1(n15598), .A2(n15599), .A3(n15600), .A4(n15601), .ZN(
        n15588) );
  NOR4_X1 U12895 ( .A1(n15590), .A2(n15591), .A3(n15592), .A4(n15593), .ZN(
        n15589) );
  OAI221_X1 U12896 ( .B1(n13480), .B2(n16532), .C1(n12776), .C2(n16526), .A(
        n15604), .ZN(n15599) );
  NAND2_X1 U12897 ( .A1(n15570), .A2(n15571), .ZN(n4903) );
  NOR4_X1 U12898 ( .A1(n15580), .A2(n15581), .A3(n15582), .A4(n15583), .ZN(
        n15570) );
  NOR4_X1 U12899 ( .A1(n15572), .A2(n15573), .A3(n15574), .A4(n15575), .ZN(
        n15571) );
  OAI221_X1 U12900 ( .B1(n13479), .B2(n16532), .C1(n12775), .C2(n16526), .A(
        n15586), .ZN(n15581) );
  NAND2_X1 U12901 ( .A1(n15552), .A2(n15553), .ZN(n4904) );
  NOR4_X1 U12902 ( .A1(n15562), .A2(n15563), .A3(n15564), .A4(n15565), .ZN(
        n15552) );
  NOR4_X1 U12903 ( .A1(n15554), .A2(n15555), .A3(n15556), .A4(n15557), .ZN(
        n15553) );
  OAI221_X1 U12904 ( .B1(n13478), .B2(n16532), .C1(n12774), .C2(n16526), .A(
        n15568), .ZN(n15563) );
  NOR2_X1 U12905 ( .A1(n12196), .A2(n12195), .ZN(n16070) );
  NOR2_X1 U12906 ( .A1(n12191), .A2(n12190), .ZN(n14862) );
  NOR3_X1 U12907 ( .A1(n12194), .A2(n12193), .A3(n12197), .ZN(n16069) );
  NOR3_X1 U12908 ( .A1(n12189), .A2(n12188), .A3(n12192), .ZN(n14861) );
  BUF_X1 U12909 ( .A(n14923), .Z(n16561) );
  BUF_X1 U12910 ( .A(n14923), .Z(n16562) );
  BUF_X1 U12911 ( .A(n14923), .Z(n16563) );
  BUF_X1 U12912 ( .A(n14923), .Z(n16564) );
  BUF_X1 U12913 ( .A(n13715), .Z(n16766) );
  BUF_X1 U12914 ( .A(n13715), .Z(n16767) );
  BUF_X1 U12915 ( .A(n13715), .Z(n16768) );
  BUF_X1 U12916 ( .A(n13715), .Z(n16769) );
  NOR2_X1 U12917 ( .A1(n16085), .A2(n16560), .ZN(n14932) );
  NOR2_X1 U12918 ( .A1(n14877), .A2(n16765), .ZN(n13720) );
  BUF_X1 U12919 ( .A(n14923), .Z(n16560) );
  BUF_X1 U12920 ( .A(n13715), .Z(n16765) );
  NAND2_X1 U12921 ( .A1(n16083), .A2(n16065), .ZN(n14925) );
  NAND2_X1 U12922 ( .A1(n14875), .A2(n14857), .ZN(n13717) );
  BUF_X1 U12923 ( .A(n16064), .Z(n16480) );
  BUF_X1 U12924 ( .A(n14856), .Z(n16685) );
  BUF_X1 U12925 ( .A(n16064), .Z(n16481) );
  BUF_X1 U12926 ( .A(n14856), .Z(n16686) );
  NAND2_X1 U12927 ( .A1(n16083), .A2(n16070), .ZN(n14919) );
  NAND2_X1 U12928 ( .A1(n14875), .A2(n14862), .ZN(n13711) );
  NAND2_X1 U12929 ( .A1(n16082), .A2(n16065), .ZN(n14924) );
  NAND2_X1 U12930 ( .A1(n14874), .A2(n14857), .ZN(n13716) );
  AND3_X1 U12931 ( .A1(n16065), .A2(n16480), .A3(n16074), .ZN(n14938) );
  AND3_X1 U12932 ( .A1(n14857), .A2(n16685), .A3(n14866), .ZN(n13730) );
  AND3_X1 U12933 ( .A1(n16066), .A2(n16069), .A3(n16480), .ZN(n14913) );
  AND3_X1 U12934 ( .A1(n14858), .A2(n14861), .A3(n16685), .ZN(n13705) );
  AND3_X1 U12935 ( .A1(n16063), .A2(n16480), .A3(n16073), .ZN(n14912) );
  AND3_X1 U12936 ( .A1(n16063), .A2(n16480), .A3(n16065), .ZN(n14898) );
  AND3_X1 U12937 ( .A1(n14855), .A2(n16685), .A3(n14865), .ZN(n13704) );
  AND3_X1 U12938 ( .A1(n14855), .A2(n16685), .A3(n14857), .ZN(n13690) );
  AND3_X1 U12939 ( .A1(n16072), .A2(n16480), .A3(n16070), .ZN(n14914) );
  AND3_X1 U12940 ( .A1(n16072), .A2(n16480), .A3(n16073), .ZN(n14902) );
  AND3_X1 U12941 ( .A1(n14864), .A2(n16685), .A3(n14862), .ZN(n13706) );
  AND3_X1 U12942 ( .A1(n14864), .A2(n16685), .A3(n14865), .ZN(n13694) );
  AND3_X1 U12943 ( .A1(n16481), .A2(n16069), .A3(n16065), .ZN(n14903) );
  AND3_X1 U12944 ( .A1(n16686), .A2(n14861), .A3(n14857), .ZN(n13695) );
  AND3_X1 U12945 ( .A1(n16481), .A2(n16066), .A3(n16067), .ZN(n14897) );
  AND3_X1 U12946 ( .A1(n16481), .A2(n16066), .A3(n16063), .ZN(n14907) );
  AND3_X1 U12947 ( .A1(n16481), .A2(n16066), .A3(n16068), .ZN(n14908) );
  AND3_X1 U12948 ( .A1(n16481), .A2(n16066), .A3(n16072), .ZN(n14937) );
  AND3_X1 U12949 ( .A1(n16481), .A2(n16066), .A3(n16074), .ZN(n14939) );
  AND3_X1 U12950 ( .A1(n16686), .A2(n14858), .A3(n14859), .ZN(n13689) );
  AND3_X1 U12951 ( .A1(n16686), .A2(n14858), .A3(n14855), .ZN(n13699) );
  AND3_X1 U12952 ( .A1(n16686), .A2(n14858), .A3(n14860), .ZN(n13700) );
  AND3_X1 U12953 ( .A1(n16686), .A2(n14858), .A3(n14864), .ZN(n13729) );
  AND3_X1 U12954 ( .A1(n16686), .A2(n14858), .A3(n14866), .ZN(n13731) );
  AND2_X1 U12955 ( .A1(n16087), .A2(n12197), .ZN(n16082) );
  AND2_X1 U12956 ( .A1(n14879), .A2(n12192), .ZN(n14874) );
  AND2_X1 U12957 ( .A1(n16083), .A2(n16066), .ZN(n14928) );
  AND2_X1 U12958 ( .A1(n16082), .A2(n16066), .ZN(n14933) );
  AND2_X1 U12959 ( .A1(n14875), .A2(n14858), .ZN(n13719) );
  AND2_X1 U12960 ( .A1(n14874), .A2(n14858), .ZN(n13724) );
  AND2_X1 U12961 ( .A1(n16083), .A2(n16073), .ZN(n14927) );
  AND2_X1 U12962 ( .A1(n16082), .A2(n16073), .ZN(n14922) );
  AND2_X1 U12963 ( .A1(n14874), .A2(n14865), .ZN(n13714) );
  AND2_X1 U12964 ( .A1(n14875), .A2(n14865), .ZN(n13725) );
  AND3_X1 U12965 ( .A1(n12194), .A2(n12193), .A3(n16480), .ZN(n16087) );
  AND3_X1 U12966 ( .A1(n12189), .A2(n12188), .A3(n16685), .ZN(n14879) );
  BUF_X1 U12967 ( .A(n13650), .Z(n17299) );
  OAI21_X1 U12968 ( .B1(n13636), .B2(n13651), .A(n17589), .ZN(n13650) );
  BUF_X1 U12969 ( .A(n13648), .Z(n17318) );
  OAI21_X1 U12970 ( .B1(n13636), .B2(n13649), .A(n17589), .ZN(n13648) );
  BUF_X1 U12971 ( .A(n13646), .Z(n17337) );
  OAI21_X1 U12972 ( .B1(n13636), .B2(n13647), .A(n17589), .ZN(n13646) );
  BUF_X1 U12973 ( .A(n13644), .Z(n17356) );
  OAI21_X1 U12974 ( .B1(n13636), .B2(n13645), .A(n17589), .ZN(n13644) );
  BUF_X1 U12975 ( .A(n13642), .Z(n17375) );
  OAI21_X1 U12976 ( .B1(n13636), .B2(n13643), .A(n17589), .ZN(n13642) );
  BUF_X1 U12977 ( .A(n13640), .Z(n17394) );
  OAI21_X1 U12978 ( .B1(n13636), .B2(n13641), .A(n17589), .ZN(n13640) );
  BUF_X1 U12979 ( .A(n13638), .Z(n17413) );
  OAI21_X1 U12980 ( .B1(n13636), .B2(n13639), .A(n17589), .ZN(n13638) );
  BUF_X1 U12981 ( .A(n13679), .Z(n16890) );
  OAI21_X1 U12982 ( .B1(n13651), .B2(n13672), .A(n17587), .ZN(n13679) );
  BUF_X1 U12983 ( .A(n13678), .Z(n16907) );
  OAI21_X1 U12984 ( .B1(n13649), .B2(n13672), .A(n17587), .ZN(n13678) );
  BUF_X1 U12985 ( .A(n13677), .Z(n16924) );
  OAI21_X1 U12986 ( .B1(n13647), .B2(n13672), .A(n17587), .ZN(n13677) );
  BUF_X1 U12987 ( .A(n13676), .Z(n16941) );
  OAI21_X1 U12988 ( .B1(n13645), .B2(n13672), .A(n17587), .ZN(n13676) );
  BUF_X1 U12989 ( .A(n13675), .Z(n16958) );
  OAI21_X1 U12990 ( .B1(n13643), .B2(n13672), .A(n17587), .ZN(n13675) );
  BUF_X1 U12991 ( .A(n13674), .Z(n16975) );
  OAI21_X1 U12992 ( .B1(n13641), .B2(n13672), .A(n17587), .ZN(n13674) );
  BUF_X1 U12993 ( .A(n13673), .Z(n16992) );
  OAI21_X1 U12994 ( .B1(n13639), .B2(n13672), .A(n17587), .ZN(n13673) );
  BUF_X1 U12995 ( .A(n13671), .Z(n17009) );
  OAI21_X1 U12996 ( .B1(n13637), .B2(n13672), .A(n17587), .ZN(n13671) );
  BUF_X1 U12997 ( .A(n13670), .Z(n17026) );
  OAI21_X1 U12998 ( .B1(n13651), .B2(n13663), .A(n17588), .ZN(n13670) );
  BUF_X1 U12999 ( .A(n13669), .Z(n17043) );
  OAI21_X1 U13000 ( .B1(n13649), .B2(n13663), .A(n17588), .ZN(n13669) );
  BUF_X1 U13001 ( .A(n13668), .Z(n17060) );
  OAI21_X1 U13002 ( .B1(n13647), .B2(n13663), .A(n17588), .ZN(n13668) );
  BUF_X1 U13003 ( .A(n13667), .Z(n17077) );
  OAI21_X1 U13004 ( .B1(n13645), .B2(n13663), .A(n17588), .ZN(n13667) );
  BUF_X1 U13005 ( .A(n13666), .Z(n17094) );
  OAI21_X1 U13006 ( .B1(n13643), .B2(n13663), .A(n17588), .ZN(n13666) );
  BUF_X1 U13007 ( .A(n13665), .Z(n17111) );
  OAI21_X1 U13008 ( .B1(n13641), .B2(n13663), .A(n17588), .ZN(n13665) );
  BUF_X1 U13009 ( .A(n13664), .Z(n17128) );
  OAI21_X1 U13010 ( .B1(n13639), .B2(n13663), .A(n17588), .ZN(n13664) );
  BUF_X1 U13011 ( .A(n13662), .Z(n17145) );
  OAI21_X1 U13012 ( .B1(n13637), .B2(n13663), .A(n17588), .ZN(n13662) );
  BUF_X1 U13013 ( .A(n13661), .Z(n17162) );
  OAI21_X1 U13014 ( .B1(n13651), .B2(n13654), .A(n17588), .ZN(n13661) );
  BUF_X1 U13015 ( .A(n13660), .Z(n17180) );
  OAI21_X1 U13016 ( .B1(n13649), .B2(n13654), .A(n17588), .ZN(n13660) );
  BUF_X1 U13017 ( .A(n13659), .Z(n17197) );
  OAI21_X1 U13018 ( .B1(n13647), .B2(n13654), .A(n17588), .ZN(n13659) );
  BUF_X1 U13019 ( .A(n13658), .Z(n17214) );
  OAI21_X1 U13020 ( .B1(n13645), .B2(n13654), .A(n17588), .ZN(n13658) );
  BUF_X1 U13021 ( .A(n13657), .Z(n17231) );
  OAI21_X1 U13022 ( .B1(n13643), .B2(n13654), .A(n17589), .ZN(n13657) );
  BUF_X1 U13023 ( .A(n13656), .Z(n17248) );
  OAI21_X1 U13024 ( .B1(n13641), .B2(n13654), .A(n17588), .ZN(n13656) );
  BUF_X1 U13025 ( .A(n13655), .Z(n17265) );
  OAI21_X1 U13026 ( .B1(n13639), .B2(n13654), .A(n17589), .ZN(n13655) );
  BUF_X1 U13027 ( .A(n13653), .Z(n17282) );
  OAI21_X1 U13028 ( .B1(n13637), .B2(n13654), .A(n17589), .ZN(n13653) );
  OAI221_X1 U13029 ( .B1(n13510), .B2(n16684), .C1(n12585), .C2(n16678), .A(
        n14982), .ZN(n14981) );
  AOI22_X1 U13030 ( .A1(n16672), .A2(n8508), .B1(n16666), .B2(n8572), .ZN(
        n14982) );
  OAI221_X1 U13031 ( .B1(n13509), .B2(n16684), .C1(n12584), .C2(n16678), .A(
        n14964), .ZN(n14963) );
  AOI22_X1 U13032 ( .A1(n16672), .A2(n8507), .B1(n16666), .B2(n8571), .ZN(
        n14964) );
  OAI221_X1 U13033 ( .B1(n13508), .B2(n16684), .C1(n12583), .C2(n16678), .A(
        n14946), .ZN(n14945) );
  AOI22_X1 U13034 ( .A1(n16672), .A2(n8506), .B1(n16666), .B2(n8570), .ZN(
        n14946) );
  OAI221_X1 U13035 ( .B1(n13507), .B2(n16684), .C1(n12582), .C2(n16678), .A(
        n14896), .ZN(n14893) );
  AOI22_X1 U13036 ( .A1(n16672), .A2(n8505), .B1(n16666), .B2(n8569), .ZN(
        n14896) );
  OAI221_X1 U13037 ( .B1(n13510), .B2(n16889), .C1(n12585), .C2(n16883), .A(
        n13774), .ZN(n13773) );
  AOI22_X1 U13038 ( .A1(n16877), .A2(n8508), .B1(n16871), .B2(n8572), .ZN(
        n13774) );
  OAI221_X1 U13039 ( .B1(n13509), .B2(n16889), .C1(n12584), .C2(n16883), .A(
        n13756), .ZN(n13755) );
  AOI22_X1 U13040 ( .A1(n16877), .A2(n8507), .B1(n16871), .B2(n8571), .ZN(
        n13756) );
  OAI221_X1 U13041 ( .B1(n13508), .B2(n16889), .C1(n12583), .C2(n16883), .A(
        n13738), .ZN(n13737) );
  AOI22_X1 U13042 ( .A1(n16877), .A2(n8506), .B1(n16871), .B2(n8570), .ZN(
        n13738) );
  OAI221_X1 U13043 ( .B1(n13507), .B2(n16889), .C1(n12582), .C2(n16883), .A(
        n13688), .ZN(n13685) );
  AOI22_X1 U13044 ( .A1(n16877), .A2(n8505), .B1(n16871), .B2(n8569), .ZN(
        n13688) );
  OAI221_X1 U13045 ( .B1(n13570), .B2(n16679), .C1(n12645), .C2(n16673), .A(
        n16062), .ZN(n16061) );
  AOI22_X1 U13046 ( .A1(n16667), .A2(n8568), .B1(n16661), .B2(n8632), .ZN(
        n16062) );
  OAI221_X1 U13047 ( .B1(n13569), .B2(n16679), .C1(n12644), .C2(n16673), .A(
        n16044), .ZN(n16043) );
  AOI22_X1 U13048 ( .A1(n16667), .A2(n8567), .B1(n16661), .B2(n8631), .ZN(
        n16044) );
  OAI221_X1 U13049 ( .B1(n13568), .B2(n16679), .C1(n12643), .C2(n16673), .A(
        n16026), .ZN(n16025) );
  AOI22_X1 U13050 ( .A1(n16667), .A2(n8566), .B1(n16661), .B2(n8630), .ZN(
        n16026) );
  OAI221_X1 U13051 ( .B1(n13567), .B2(n16679), .C1(n12642), .C2(n16673), .A(
        n16008), .ZN(n16007) );
  AOI22_X1 U13052 ( .A1(n16667), .A2(n8565), .B1(n16661), .B2(n8629), .ZN(
        n16008) );
  OAI221_X1 U13053 ( .B1(n13566), .B2(n16679), .C1(n12641), .C2(n16673), .A(
        n15990), .ZN(n15989) );
  AOI22_X1 U13054 ( .A1(n16667), .A2(n8564), .B1(n16661), .B2(n8628), .ZN(
        n15990) );
  OAI221_X1 U13055 ( .B1(n13565), .B2(n16679), .C1(n12640), .C2(n16673), .A(
        n15972), .ZN(n15971) );
  AOI22_X1 U13056 ( .A1(n16667), .A2(n8563), .B1(n16661), .B2(n8627), .ZN(
        n15972) );
  OAI221_X1 U13057 ( .B1(n13564), .B2(n16679), .C1(n12639), .C2(n16673), .A(
        n15954), .ZN(n15953) );
  AOI22_X1 U13058 ( .A1(n16667), .A2(n8562), .B1(n16661), .B2(n8626), .ZN(
        n15954) );
  OAI221_X1 U13059 ( .B1(n13563), .B2(n16679), .C1(n12638), .C2(n16673), .A(
        n15936), .ZN(n15935) );
  AOI22_X1 U13060 ( .A1(n16667), .A2(n8561), .B1(n16661), .B2(n8625), .ZN(
        n15936) );
  OAI221_X1 U13061 ( .B1(n13562), .B2(n16679), .C1(n12637), .C2(n16673), .A(
        n15918), .ZN(n15917) );
  AOI22_X1 U13062 ( .A1(n16667), .A2(n8560), .B1(n16661), .B2(n8624), .ZN(
        n15918) );
  OAI221_X1 U13063 ( .B1(n13561), .B2(n16679), .C1(n12636), .C2(n16673), .A(
        n15900), .ZN(n15899) );
  AOI22_X1 U13064 ( .A1(n16667), .A2(n8559), .B1(n16661), .B2(n8623), .ZN(
        n15900) );
  OAI221_X1 U13065 ( .B1(n13560), .B2(n16679), .C1(n12635), .C2(n16673), .A(
        n15882), .ZN(n15881) );
  AOI22_X1 U13066 ( .A1(n16667), .A2(n8558), .B1(n16661), .B2(n8622), .ZN(
        n15882) );
  OAI221_X1 U13067 ( .B1(n13559), .B2(n16679), .C1(n12634), .C2(n16673), .A(
        n15864), .ZN(n15863) );
  AOI22_X1 U13068 ( .A1(n16667), .A2(n8557), .B1(n16661), .B2(n8621), .ZN(
        n15864) );
  OAI221_X1 U13069 ( .B1(n13558), .B2(n16680), .C1(n12633), .C2(n16674), .A(
        n15846), .ZN(n15845) );
  AOI22_X1 U13070 ( .A1(n16668), .A2(n8556), .B1(n16662), .B2(n8620), .ZN(
        n15846) );
  OAI221_X1 U13071 ( .B1(n13557), .B2(n16680), .C1(n12632), .C2(n16674), .A(
        n15828), .ZN(n15827) );
  AOI22_X1 U13072 ( .A1(n16668), .A2(n8555), .B1(n16662), .B2(n8619), .ZN(
        n15828) );
  OAI221_X1 U13073 ( .B1(n13556), .B2(n16680), .C1(n12631), .C2(n16674), .A(
        n15810), .ZN(n15809) );
  AOI22_X1 U13074 ( .A1(n16668), .A2(n8554), .B1(n16662), .B2(n8618), .ZN(
        n15810) );
  OAI221_X1 U13075 ( .B1(n13555), .B2(n16680), .C1(n12630), .C2(n16674), .A(
        n15792), .ZN(n15791) );
  AOI22_X1 U13076 ( .A1(n16668), .A2(n8553), .B1(n16662), .B2(n8617), .ZN(
        n15792) );
  OAI221_X1 U13077 ( .B1(n13554), .B2(n16680), .C1(n12629), .C2(n16674), .A(
        n15774), .ZN(n15773) );
  AOI22_X1 U13078 ( .A1(n16668), .A2(n8552), .B1(n16662), .B2(n8616), .ZN(
        n15774) );
  OAI221_X1 U13079 ( .B1(n13553), .B2(n16680), .C1(n12628), .C2(n16674), .A(
        n15756), .ZN(n15755) );
  AOI22_X1 U13080 ( .A1(n16668), .A2(n8551), .B1(n16662), .B2(n8615), .ZN(
        n15756) );
  OAI221_X1 U13081 ( .B1(n13552), .B2(n16680), .C1(n12627), .C2(n16674), .A(
        n15738), .ZN(n15737) );
  AOI22_X1 U13082 ( .A1(n16668), .A2(n8550), .B1(n16662), .B2(n8614), .ZN(
        n15738) );
  OAI221_X1 U13083 ( .B1(n13551), .B2(n16680), .C1(n12626), .C2(n16674), .A(
        n15720), .ZN(n15719) );
  AOI22_X1 U13084 ( .A1(n16668), .A2(n8549), .B1(n16662), .B2(n8613), .ZN(
        n15720) );
  OAI221_X1 U13085 ( .B1(n13550), .B2(n16680), .C1(n12625), .C2(n16674), .A(
        n15702), .ZN(n15701) );
  AOI22_X1 U13086 ( .A1(n16668), .A2(n8548), .B1(n16662), .B2(n8612), .ZN(
        n15702) );
  OAI221_X1 U13087 ( .B1(n13549), .B2(n16680), .C1(n12624), .C2(n16674), .A(
        n15684), .ZN(n15683) );
  AOI22_X1 U13088 ( .A1(n16668), .A2(n8547), .B1(n16662), .B2(n8611), .ZN(
        n15684) );
  OAI221_X1 U13089 ( .B1(n13548), .B2(n16680), .C1(n12623), .C2(n16674), .A(
        n15666), .ZN(n15665) );
  AOI22_X1 U13090 ( .A1(n16668), .A2(n8546), .B1(n16662), .B2(n8610), .ZN(
        n15666) );
  OAI221_X1 U13091 ( .B1(n13547), .B2(n16680), .C1(n12622), .C2(n16674), .A(
        n15648), .ZN(n15647) );
  AOI22_X1 U13092 ( .A1(n16668), .A2(n8545), .B1(n16662), .B2(n8609), .ZN(
        n15648) );
  OAI221_X1 U13093 ( .B1(n13546), .B2(n16681), .C1(n12621), .C2(n16675), .A(
        n15630), .ZN(n15629) );
  AOI22_X1 U13094 ( .A1(n16669), .A2(n8544), .B1(n16663), .B2(n8608), .ZN(
        n15630) );
  OAI221_X1 U13095 ( .B1(n13545), .B2(n16681), .C1(n12620), .C2(n16675), .A(
        n15612), .ZN(n15611) );
  AOI22_X1 U13096 ( .A1(n16669), .A2(n8543), .B1(n16663), .B2(n8607), .ZN(
        n15612) );
  OAI221_X1 U13097 ( .B1(n13544), .B2(n16681), .C1(n12619), .C2(n16675), .A(
        n15594), .ZN(n15593) );
  AOI22_X1 U13098 ( .A1(n16669), .A2(n8542), .B1(n16663), .B2(n8606), .ZN(
        n15594) );
  OAI221_X1 U13099 ( .B1(n13543), .B2(n16681), .C1(n12618), .C2(n16675), .A(
        n15576), .ZN(n15575) );
  AOI22_X1 U13100 ( .A1(n16669), .A2(n8541), .B1(n16663), .B2(n8605), .ZN(
        n15576) );
  OAI221_X1 U13101 ( .B1(n13542), .B2(n16681), .C1(n12617), .C2(n16675), .A(
        n15558), .ZN(n15557) );
  AOI22_X1 U13102 ( .A1(n16669), .A2(n8540), .B1(n16663), .B2(n8604), .ZN(
        n15558) );
  OAI221_X1 U13103 ( .B1(n13541), .B2(n16681), .C1(n12616), .C2(n16675), .A(
        n15540), .ZN(n15539) );
  AOI22_X1 U13104 ( .A1(n16669), .A2(n8539), .B1(n16663), .B2(n8603), .ZN(
        n15540) );
  OAI221_X1 U13105 ( .B1(n13540), .B2(n16681), .C1(n12615), .C2(n16675), .A(
        n15522), .ZN(n15521) );
  AOI22_X1 U13106 ( .A1(n16669), .A2(n8538), .B1(n16663), .B2(n8602), .ZN(
        n15522) );
  OAI221_X1 U13107 ( .B1(n13539), .B2(n16681), .C1(n12614), .C2(n16675), .A(
        n15504), .ZN(n15503) );
  AOI22_X1 U13108 ( .A1(n16669), .A2(n8537), .B1(n16663), .B2(n8601), .ZN(
        n15504) );
  OAI221_X1 U13109 ( .B1(n13538), .B2(n16681), .C1(n12613), .C2(n16675), .A(
        n15486), .ZN(n15485) );
  AOI22_X1 U13110 ( .A1(n16669), .A2(n8536), .B1(n16663), .B2(n8600), .ZN(
        n15486) );
  OAI221_X1 U13111 ( .B1(n13537), .B2(n16681), .C1(n12612), .C2(n16675), .A(
        n15468), .ZN(n15467) );
  AOI22_X1 U13112 ( .A1(n16669), .A2(n8535), .B1(n16663), .B2(n8599), .ZN(
        n15468) );
  OAI221_X1 U13113 ( .B1(n13536), .B2(n16681), .C1(n12611), .C2(n16675), .A(
        n15450), .ZN(n15449) );
  AOI22_X1 U13114 ( .A1(n16669), .A2(n8534), .B1(n16663), .B2(n8598), .ZN(
        n15450) );
  OAI221_X1 U13115 ( .B1(n13535), .B2(n16681), .C1(n12610), .C2(n16675), .A(
        n15432), .ZN(n15431) );
  AOI22_X1 U13116 ( .A1(n16669), .A2(n8533), .B1(n16663), .B2(n8597), .ZN(
        n15432) );
  OAI221_X1 U13117 ( .B1(n13534), .B2(n16682), .C1(n12609), .C2(n16676), .A(
        n15414), .ZN(n15413) );
  AOI22_X1 U13118 ( .A1(n16670), .A2(n8532), .B1(n16664), .B2(n8596), .ZN(
        n15414) );
  OAI221_X1 U13119 ( .B1(n13533), .B2(n16682), .C1(n12608), .C2(n16676), .A(
        n15396), .ZN(n15395) );
  AOI22_X1 U13120 ( .A1(n16670), .A2(n8531), .B1(n16664), .B2(n8595), .ZN(
        n15396) );
  OAI221_X1 U13121 ( .B1(n13532), .B2(n16682), .C1(n12607), .C2(n16676), .A(
        n15378), .ZN(n15377) );
  AOI22_X1 U13122 ( .A1(n16670), .A2(n8530), .B1(n16664), .B2(n8594), .ZN(
        n15378) );
  OAI221_X1 U13123 ( .B1(n13531), .B2(n16682), .C1(n12606), .C2(n16676), .A(
        n15360), .ZN(n15359) );
  AOI22_X1 U13124 ( .A1(n16670), .A2(n8529), .B1(n16664), .B2(n8593), .ZN(
        n15360) );
  OAI221_X1 U13125 ( .B1(n13530), .B2(n16682), .C1(n12605), .C2(n16676), .A(
        n15342), .ZN(n15341) );
  AOI22_X1 U13126 ( .A1(n16670), .A2(n8528), .B1(n16664), .B2(n8592), .ZN(
        n15342) );
  OAI221_X1 U13127 ( .B1(n13529), .B2(n16682), .C1(n12604), .C2(n16676), .A(
        n15324), .ZN(n15323) );
  AOI22_X1 U13128 ( .A1(n16670), .A2(n8527), .B1(n16664), .B2(n8591), .ZN(
        n15324) );
  OAI221_X1 U13129 ( .B1(n13528), .B2(n16682), .C1(n12603), .C2(n16676), .A(
        n15306), .ZN(n15305) );
  AOI22_X1 U13130 ( .A1(n16670), .A2(n8526), .B1(n16664), .B2(n8590), .ZN(
        n15306) );
  OAI221_X1 U13131 ( .B1(n13527), .B2(n16682), .C1(n12602), .C2(n16676), .A(
        n15288), .ZN(n15287) );
  AOI22_X1 U13132 ( .A1(n16670), .A2(n8525), .B1(n16664), .B2(n8589), .ZN(
        n15288) );
  OAI221_X1 U13133 ( .B1(n13526), .B2(n16682), .C1(n12601), .C2(n16676), .A(
        n15270), .ZN(n15269) );
  AOI22_X1 U13134 ( .A1(n16670), .A2(n8524), .B1(n16664), .B2(n8588), .ZN(
        n15270) );
  OAI221_X1 U13135 ( .B1(n13525), .B2(n16682), .C1(n12600), .C2(n16676), .A(
        n15252), .ZN(n15251) );
  AOI22_X1 U13136 ( .A1(n16670), .A2(n8523), .B1(n16664), .B2(n8587), .ZN(
        n15252) );
  OAI221_X1 U13137 ( .B1(n13524), .B2(n16682), .C1(n12599), .C2(n16676), .A(
        n15234), .ZN(n15233) );
  AOI22_X1 U13138 ( .A1(n16670), .A2(n8522), .B1(n16664), .B2(n8586), .ZN(
        n15234) );
  OAI221_X1 U13139 ( .B1(n13523), .B2(n16682), .C1(n12598), .C2(n16676), .A(
        n15216), .ZN(n15215) );
  AOI22_X1 U13140 ( .A1(n16670), .A2(n8521), .B1(n16664), .B2(n8585), .ZN(
        n15216) );
  OAI221_X1 U13141 ( .B1(n13570), .B2(n16884), .C1(n12645), .C2(n16878), .A(
        n14854), .ZN(n14853) );
  AOI22_X1 U13142 ( .A1(n16872), .A2(n8568), .B1(n16866), .B2(n8632), .ZN(
        n14854) );
  OAI221_X1 U13143 ( .B1(n13569), .B2(n16884), .C1(n12644), .C2(n16878), .A(
        n14836), .ZN(n14835) );
  AOI22_X1 U13144 ( .A1(n16872), .A2(n8567), .B1(n16866), .B2(n8631), .ZN(
        n14836) );
  OAI221_X1 U13145 ( .B1(n13568), .B2(n16884), .C1(n12643), .C2(n16878), .A(
        n14818), .ZN(n14817) );
  AOI22_X1 U13146 ( .A1(n16872), .A2(n8566), .B1(n16866), .B2(n8630), .ZN(
        n14818) );
  OAI221_X1 U13147 ( .B1(n13567), .B2(n16884), .C1(n12642), .C2(n16878), .A(
        n14800), .ZN(n14799) );
  AOI22_X1 U13148 ( .A1(n16872), .A2(n8565), .B1(n16866), .B2(n8629), .ZN(
        n14800) );
  OAI221_X1 U13149 ( .B1(n13566), .B2(n16884), .C1(n12641), .C2(n16878), .A(
        n14782), .ZN(n14781) );
  AOI22_X1 U13150 ( .A1(n16872), .A2(n8564), .B1(n16866), .B2(n8628), .ZN(
        n14782) );
  OAI221_X1 U13151 ( .B1(n13565), .B2(n16884), .C1(n12640), .C2(n16878), .A(
        n14764), .ZN(n14763) );
  AOI22_X1 U13152 ( .A1(n16872), .A2(n8563), .B1(n16866), .B2(n8627), .ZN(
        n14764) );
  OAI221_X1 U13153 ( .B1(n13564), .B2(n16884), .C1(n12639), .C2(n16878), .A(
        n14746), .ZN(n14745) );
  AOI22_X1 U13154 ( .A1(n16872), .A2(n8562), .B1(n16866), .B2(n8626), .ZN(
        n14746) );
  OAI221_X1 U13155 ( .B1(n13563), .B2(n16884), .C1(n12638), .C2(n16878), .A(
        n14728), .ZN(n14727) );
  AOI22_X1 U13156 ( .A1(n16872), .A2(n8561), .B1(n16866), .B2(n8625), .ZN(
        n14728) );
  OAI221_X1 U13157 ( .B1(n13562), .B2(n16884), .C1(n12637), .C2(n16878), .A(
        n14710), .ZN(n14709) );
  AOI22_X1 U13158 ( .A1(n16872), .A2(n8560), .B1(n16866), .B2(n8624), .ZN(
        n14710) );
  OAI221_X1 U13159 ( .B1(n13561), .B2(n16884), .C1(n12636), .C2(n16878), .A(
        n14692), .ZN(n14691) );
  AOI22_X1 U13160 ( .A1(n16872), .A2(n8559), .B1(n16866), .B2(n8623), .ZN(
        n14692) );
  OAI221_X1 U13161 ( .B1(n13560), .B2(n16884), .C1(n12635), .C2(n16878), .A(
        n14674), .ZN(n14673) );
  AOI22_X1 U13162 ( .A1(n16872), .A2(n8558), .B1(n16866), .B2(n8622), .ZN(
        n14674) );
  OAI221_X1 U13163 ( .B1(n13559), .B2(n16884), .C1(n12634), .C2(n16878), .A(
        n14656), .ZN(n14655) );
  AOI22_X1 U13164 ( .A1(n16872), .A2(n8557), .B1(n16866), .B2(n8621), .ZN(
        n14656) );
  OAI221_X1 U13165 ( .B1(n13558), .B2(n16885), .C1(n12633), .C2(n16879), .A(
        n14638), .ZN(n14637) );
  AOI22_X1 U13166 ( .A1(n16873), .A2(n8556), .B1(n16867), .B2(n8620), .ZN(
        n14638) );
  OAI221_X1 U13167 ( .B1(n13557), .B2(n16885), .C1(n12632), .C2(n16879), .A(
        n14620), .ZN(n14619) );
  AOI22_X1 U13168 ( .A1(n16873), .A2(n8555), .B1(n16867), .B2(n8619), .ZN(
        n14620) );
  OAI221_X1 U13169 ( .B1(n13556), .B2(n16885), .C1(n12631), .C2(n16879), .A(
        n14602), .ZN(n14601) );
  AOI22_X1 U13170 ( .A1(n16873), .A2(n8554), .B1(n16867), .B2(n8618), .ZN(
        n14602) );
  OAI221_X1 U13171 ( .B1(n13555), .B2(n16885), .C1(n12630), .C2(n16879), .A(
        n14584), .ZN(n14583) );
  AOI22_X1 U13172 ( .A1(n16873), .A2(n8553), .B1(n16867), .B2(n8617), .ZN(
        n14584) );
  OAI221_X1 U13173 ( .B1(n13554), .B2(n16885), .C1(n12629), .C2(n16879), .A(
        n14566), .ZN(n14565) );
  AOI22_X1 U13174 ( .A1(n16873), .A2(n8552), .B1(n16867), .B2(n8616), .ZN(
        n14566) );
  OAI221_X1 U13175 ( .B1(n13553), .B2(n16885), .C1(n12628), .C2(n16879), .A(
        n14548), .ZN(n14547) );
  AOI22_X1 U13176 ( .A1(n16873), .A2(n8551), .B1(n16867), .B2(n8615), .ZN(
        n14548) );
  OAI221_X1 U13177 ( .B1(n13552), .B2(n16885), .C1(n12627), .C2(n16879), .A(
        n14530), .ZN(n14529) );
  AOI22_X1 U13178 ( .A1(n16873), .A2(n8550), .B1(n16867), .B2(n8614), .ZN(
        n14530) );
  OAI221_X1 U13179 ( .B1(n13551), .B2(n16885), .C1(n12626), .C2(n16879), .A(
        n14512), .ZN(n14511) );
  AOI22_X1 U13180 ( .A1(n16873), .A2(n8549), .B1(n16867), .B2(n8613), .ZN(
        n14512) );
  OAI221_X1 U13181 ( .B1(n13550), .B2(n16885), .C1(n12625), .C2(n16879), .A(
        n14494), .ZN(n14493) );
  AOI22_X1 U13182 ( .A1(n16873), .A2(n8548), .B1(n16867), .B2(n8612), .ZN(
        n14494) );
  OAI221_X1 U13183 ( .B1(n13549), .B2(n16885), .C1(n12624), .C2(n16879), .A(
        n14476), .ZN(n14475) );
  AOI22_X1 U13184 ( .A1(n16873), .A2(n8547), .B1(n16867), .B2(n8611), .ZN(
        n14476) );
  OAI221_X1 U13185 ( .B1(n13548), .B2(n16885), .C1(n12623), .C2(n16879), .A(
        n14458), .ZN(n14457) );
  AOI22_X1 U13186 ( .A1(n16873), .A2(n8546), .B1(n16867), .B2(n8610), .ZN(
        n14458) );
  OAI221_X1 U13187 ( .B1(n13547), .B2(n16885), .C1(n12622), .C2(n16879), .A(
        n14440), .ZN(n14439) );
  AOI22_X1 U13188 ( .A1(n16873), .A2(n8545), .B1(n16867), .B2(n8609), .ZN(
        n14440) );
  OAI221_X1 U13189 ( .B1(n13546), .B2(n16886), .C1(n12621), .C2(n16880), .A(
        n14422), .ZN(n14421) );
  AOI22_X1 U13190 ( .A1(n16874), .A2(n8544), .B1(n16868), .B2(n8608), .ZN(
        n14422) );
  OAI221_X1 U13191 ( .B1(n13545), .B2(n16886), .C1(n12620), .C2(n16880), .A(
        n14404), .ZN(n14403) );
  AOI22_X1 U13192 ( .A1(n16874), .A2(n8543), .B1(n16868), .B2(n8607), .ZN(
        n14404) );
  OAI221_X1 U13193 ( .B1(n13544), .B2(n16886), .C1(n12619), .C2(n16880), .A(
        n14386), .ZN(n14385) );
  AOI22_X1 U13194 ( .A1(n16874), .A2(n8542), .B1(n16868), .B2(n8606), .ZN(
        n14386) );
  OAI221_X1 U13195 ( .B1(n13543), .B2(n16886), .C1(n12618), .C2(n16880), .A(
        n14368), .ZN(n14367) );
  AOI22_X1 U13196 ( .A1(n16874), .A2(n8541), .B1(n16868), .B2(n8605), .ZN(
        n14368) );
  OAI221_X1 U13197 ( .B1(n13542), .B2(n16886), .C1(n12617), .C2(n16880), .A(
        n14350), .ZN(n14349) );
  AOI22_X1 U13198 ( .A1(n16874), .A2(n8540), .B1(n16868), .B2(n8604), .ZN(
        n14350) );
  OAI221_X1 U13199 ( .B1(n13541), .B2(n16886), .C1(n12616), .C2(n16880), .A(
        n14332), .ZN(n14331) );
  AOI22_X1 U13200 ( .A1(n16874), .A2(n8539), .B1(n16868), .B2(n8603), .ZN(
        n14332) );
  OAI221_X1 U13201 ( .B1(n13540), .B2(n16886), .C1(n12615), .C2(n16880), .A(
        n14314), .ZN(n14313) );
  AOI22_X1 U13202 ( .A1(n16874), .A2(n8538), .B1(n16868), .B2(n8602), .ZN(
        n14314) );
  OAI221_X1 U13203 ( .B1(n13539), .B2(n16886), .C1(n12614), .C2(n16880), .A(
        n14296), .ZN(n14295) );
  AOI22_X1 U13204 ( .A1(n16874), .A2(n8537), .B1(n16868), .B2(n8601), .ZN(
        n14296) );
  OAI221_X1 U13205 ( .B1(n13538), .B2(n16886), .C1(n12613), .C2(n16880), .A(
        n14278), .ZN(n14277) );
  AOI22_X1 U13206 ( .A1(n16874), .A2(n8536), .B1(n16868), .B2(n8600), .ZN(
        n14278) );
  OAI221_X1 U13207 ( .B1(n13537), .B2(n16886), .C1(n12612), .C2(n16880), .A(
        n14260), .ZN(n14259) );
  AOI22_X1 U13208 ( .A1(n16874), .A2(n8535), .B1(n16868), .B2(n8599), .ZN(
        n14260) );
  OAI221_X1 U13209 ( .B1(n13536), .B2(n16886), .C1(n12611), .C2(n16880), .A(
        n14242), .ZN(n14241) );
  AOI22_X1 U13210 ( .A1(n16874), .A2(n8534), .B1(n16868), .B2(n8598), .ZN(
        n14242) );
  OAI221_X1 U13211 ( .B1(n13535), .B2(n16886), .C1(n12610), .C2(n16880), .A(
        n14224), .ZN(n14223) );
  AOI22_X1 U13212 ( .A1(n16874), .A2(n8533), .B1(n16868), .B2(n8597), .ZN(
        n14224) );
  OAI221_X1 U13213 ( .B1(n13534), .B2(n16887), .C1(n12609), .C2(n16881), .A(
        n14206), .ZN(n14205) );
  AOI22_X1 U13214 ( .A1(n16875), .A2(n8532), .B1(n16869), .B2(n8596), .ZN(
        n14206) );
  OAI221_X1 U13215 ( .B1(n13533), .B2(n16887), .C1(n12608), .C2(n16881), .A(
        n14188), .ZN(n14187) );
  AOI22_X1 U13216 ( .A1(n16875), .A2(n8531), .B1(n16869), .B2(n8595), .ZN(
        n14188) );
  OAI221_X1 U13217 ( .B1(n13532), .B2(n16887), .C1(n12607), .C2(n16881), .A(
        n14170), .ZN(n14169) );
  AOI22_X1 U13218 ( .A1(n16875), .A2(n8530), .B1(n16869), .B2(n8594), .ZN(
        n14170) );
  OAI221_X1 U13219 ( .B1(n13531), .B2(n16887), .C1(n12606), .C2(n16881), .A(
        n14152), .ZN(n14151) );
  AOI22_X1 U13220 ( .A1(n16875), .A2(n8529), .B1(n16869), .B2(n8593), .ZN(
        n14152) );
  OAI221_X1 U13221 ( .B1(n13530), .B2(n16887), .C1(n12605), .C2(n16881), .A(
        n14134), .ZN(n14133) );
  AOI22_X1 U13222 ( .A1(n16875), .A2(n8528), .B1(n16869), .B2(n8592), .ZN(
        n14134) );
  OAI221_X1 U13223 ( .B1(n13529), .B2(n16887), .C1(n12604), .C2(n16881), .A(
        n14116), .ZN(n14115) );
  AOI22_X1 U13224 ( .A1(n16875), .A2(n8527), .B1(n16869), .B2(n8591), .ZN(
        n14116) );
  OAI221_X1 U13225 ( .B1(n13528), .B2(n16887), .C1(n12603), .C2(n16881), .A(
        n14098), .ZN(n14097) );
  AOI22_X1 U13226 ( .A1(n16875), .A2(n8526), .B1(n16869), .B2(n8590), .ZN(
        n14098) );
  OAI221_X1 U13227 ( .B1(n13527), .B2(n16887), .C1(n12602), .C2(n16881), .A(
        n14080), .ZN(n14079) );
  AOI22_X1 U13228 ( .A1(n16875), .A2(n8525), .B1(n16869), .B2(n8589), .ZN(
        n14080) );
  OAI221_X1 U13229 ( .B1(n13526), .B2(n16887), .C1(n12601), .C2(n16881), .A(
        n14062), .ZN(n14061) );
  AOI22_X1 U13230 ( .A1(n16875), .A2(n8524), .B1(n16869), .B2(n8588), .ZN(
        n14062) );
  OAI221_X1 U13231 ( .B1(n13525), .B2(n16887), .C1(n12600), .C2(n16881), .A(
        n14044), .ZN(n14043) );
  AOI22_X1 U13232 ( .A1(n16875), .A2(n8523), .B1(n16869), .B2(n8587), .ZN(
        n14044) );
  OAI221_X1 U13233 ( .B1(n13524), .B2(n16887), .C1(n12599), .C2(n16881), .A(
        n14026), .ZN(n14025) );
  AOI22_X1 U13234 ( .A1(n16875), .A2(n8522), .B1(n16869), .B2(n8586), .ZN(
        n14026) );
  OAI221_X1 U13235 ( .B1(n13523), .B2(n16887), .C1(n12598), .C2(n16881), .A(
        n14008), .ZN(n14007) );
  AOI22_X1 U13236 ( .A1(n16875), .A2(n8521), .B1(n16869), .B2(n8585), .ZN(
        n14008) );
  OAI221_X1 U13237 ( .B1(n13522), .B2(n16683), .C1(n12597), .C2(n16677), .A(
        n15198), .ZN(n15197) );
  AOI22_X1 U13238 ( .A1(n16671), .A2(n8520), .B1(n16665), .B2(n8584), .ZN(
        n15198) );
  OAI221_X1 U13239 ( .B1(n13521), .B2(n16683), .C1(n12596), .C2(n16677), .A(
        n15180), .ZN(n15179) );
  AOI22_X1 U13240 ( .A1(n16671), .A2(n8519), .B1(n16665), .B2(n8583), .ZN(
        n15180) );
  OAI221_X1 U13241 ( .B1(n13520), .B2(n16683), .C1(n12595), .C2(n16677), .A(
        n15162), .ZN(n15161) );
  AOI22_X1 U13242 ( .A1(n16671), .A2(n8518), .B1(n16665), .B2(n8582), .ZN(
        n15162) );
  OAI221_X1 U13243 ( .B1(n13519), .B2(n16683), .C1(n12594), .C2(n16677), .A(
        n15144), .ZN(n15143) );
  AOI22_X1 U13244 ( .A1(n16671), .A2(n8517), .B1(n16665), .B2(n8581), .ZN(
        n15144) );
  OAI221_X1 U13245 ( .B1(n13518), .B2(n16683), .C1(n12593), .C2(n16677), .A(
        n15126), .ZN(n15125) );
  AOI22_X1 U13246 ( .A1(n16671), .A2(n8516), .B1(n16665), .B2(n8580), .ZN(
        n15126) );
  OAI221_X1 U13247 ( .B1(n13517), .B2(n16683), .C1(n12592), .C2(n16677), .A(
        n15108), .ZN(n15107) );
  AOI22_X1 U13248 ( .A1(n16671), .A2(n8515), .B1(n16665), .B2(n8579), .ZN(
        n15108) );
  OAI221_X1 U13249 ( .B1(n13516), .B2(n16683), .C1(n12591), .C2(n16677), .A(
        n15090), .ZN(n15089) );
  AOI22_X1 U13250 ( .A1(n16671), .A2(n8514), .B1(n16665), .B2(n8578), .ZN(
        n15090) );
  OAI221_X1 U13251 ( .B1(n13515), .B2(n16683), .C1(n12590), .C2(n16677), .A(
        n15072), .ZN(n15071) );
  AOI22_X1 U13252 ( .A1(n16671), .A2(n8513), .B1(n16665), .B2(n8577), .ZN(
        n15072) );
  OAI221_X1 U13253 ( .B1(n13514), .B2(n16683), .C1(n12589), .C2(n16677), .A(
        n15054), .ZN(n15053) );
  AOI22_X1 U13254 ( .A1(n16671), .A2(n8512), .B1(n16665), .B2(n8576), .ZN(
        n15054) );
  OAI221_X1 U13255 ( .B1(n13513), .B2(n16683), .C1(n12588), .C2(n16677), .A(
        n15036), .ZN(n15035) );
  AOI22_X1 U13256 ( .A1(n16671), .A2(n8511), .B1(n16665), .B2(n8575), .ZN(
        n15036) );
  OAI221_X1 U13257 ( .B1(n13512), .B2(n16683), .C1(n12587), .C2(n16677), .A(
        n15018), .ZN(n15017) );
  AOI22_X1 U13258 ( .A1(n16671), .A2(n8510), .B1(n16665), .B2(n8574), .ZN(
        n15018) );
  OAI221_X1 U13259 ( .B1(n13511), .B2(n16683), .C1(n12586), .C2(n16677), .A(
        n15000), .ZN(n14999) );
  AOI22_X1 U13260 ( .A1(n16671), .A2(n8509), .B1(n16665), .B2(n8573), .ZN(
        n15000) );
  OAI221_X1 U13261 ( .B1(n13522), .B2(n16888), .C1(n12597), .C2(n16882), .A(
        n13990), .ZN(n13989) );
  AOI22_X1 U13262 ( .A1(n16876), .A2(n8520), .B1(n16870), .B2(n8584), .ZN(
        n13990) );
  OAI221_X1 U13263 ( .B1(n13521), .B2(n16888), .C1(n12596), .C2(n16882), .A(
        n13972), .ZN(n13971) );
  AOI22_X1 U13264 ( .A1(n16876), .A2(n8519), .B1(n16870), .B2(n8583), .ZN(
        n13972) );
  OAI221_X1 U13265 ( .B1(n13520), .B2(n16888), .C1(n12595), .C2(n16882), .A(
        n13954), .ZN(n13953) );
  AOI22_X1 U13266 ( .A1(n16876), .A2(n8518), .B1(n16870), .B2(n8582), .ZN(
        n13954) );
  OAI221_X1 U13267 ( .B1(n13519), .B2(n16888), .C1(n12594), .C2(n16882), .A(
        n13936), .ZN(n13935) );
  AOI22_X1 U13268 ( .A1(n16876), .A2(n8517), .B1(n16870), .B2(n8581), .ZN(
        n13936) );
  OAI221_X1 U13269 ( .B1(n13518), .B2(n16888), .C1(n12593), .C2(n16882), .A(
        n13918), .ZN(n13917) );
  AOI22_X1 U13270 ( .A1(n16876), .A2(n8516), .B1(n16870), .B2(n8580), .ZN(
        n13918) );
  OAI221_X1 U13271 ( .B1(n13517), .B2(n16888), .C1(n12592), .C2(n16882), .A(
        n13900), .ZN(n13899) );
  AOI22_X1 U13272 ( .A1(n16876), .A2(n8515), .B1(n16870), .B2(n8579), .ZN(
        n13900) );
  OAI221_X1 U13273 ( .B1(n13516), .B2(n16888), .C1(n12591), .C2(n16882), .A(
        n13882), .ZN(n13881) );
  AOI22_X1 U13274 ( .A1(n16876), .A2(n8514), .B1(n16870), .B2(n8578), .ZN(
        n13882) );
  OAI221_X1 U13275 ( .B1(n13515), .B2(n16888), .C1(n12590), .C2(n16882), .A(
        n13864), .ZN(n13863) );
  AOI22_X1 U13276 ( .A1(n16876), .A2(n8513), .B1(n16870), .B2(n8577), .ZN(
        n13864) );
  OAI221_X1 U13277 ( .B1(n13514), .B2(n16888), .C1(n12589), .C2(n16882), .A(
        n13846), .ZN(n13845) );
  AOI22_X1 U13278 ( .A1(n16876), .A2(n8512), .B1(n16870), .B2(n8576), .ZN(
        n13846) );
  OAI221_X1 U13279 ( .B1(n13513), .B2(n16888), .C1(n12588), .C2(n16882), .A(
        n13828), .ZN(n13827) );
  AOI22_X1 U13280 ( .A1(n16876), .A2(n8511), .B1(n16870), .B2(n8575), .ZN(
        n13828) );
  OAI221_X1 U13281 ( .B1(n13512), .B2(n16888), .C1(n12587), .C2(n16882), .A(
        n13810), .ZN(n13809) );
  AOI22_X1 U13282 ( .A1(n16876), .A2(n8510), .B1(n16870), .B2(n8574), .ZN(
        n13810) );
  OAI221_X1 U13283 ( .B1(n13511), .B2(n16888), .C1(n12586), .C2(n16882), .A(
        n13792), .ZN(n13791) );
  AOI22_X1 U13284 ( .A1(n16876), .A2(n8509), .B1(n16870), .B2(n8573), .ZN(
        n13792) );
  OAI221_X1 U13285 ( .B1(n16351), .B2(n16555), .C1(n16352), .C2(n16549), .A(
        n15855), .ZN(n15852) );
  AOI22_X1 U13286 ( .A1(n16546), .A2(n12441), .B1(n16537), .B2(n12313), .ZN(
        n15855) );
  OAI221_X1 U13287 ( .B1(n16346), .B2(n16555), .C1(n16347), .C2(n16549), .A(
        n15837), .ZN(n15834) );
  AOI22_X1 U13288 ( .A1(n16546), .A2(n12440), .B1(n16537), .B2(n12312), .ZN(
        n15837) );
  OAI221_X1 U13289 ( .B1(n16341), .B2(n16555), .C1(n16342), .C2(n16549), .A(
        n15819), .ZN(n15816) );
  AOI22_X1 U13290 ( .A1(n16546), .A2(n12439), .B1(n16537), .B2(n12311), .ZN(
        n15819) );
  OAI221_X1 U13291 ( .B1(n16336), .B2(n16555), .C1(n16337), .C2(n16549), .A(
        n15801), .ZN(n15798) );
  AOI22_X1 U13292 ( .A1(n16546), .A2(n12438), .B1(n16537), .B2(n12310), .ZN(
        n15801) );
  OAI221_X1 U13293 ( .B1(n16331), .B2(n16555), .C1(n16332), .C2(n16549), .A(
        n15783), .ZN(n15780) );
  AOI22_X1 U13294 ( .A1(n16545), .A2(n12437), .B1(n16537), .B2(n12309), .ZN(
        n15783) );
  OAI221_X1 U13295 ( .B1(n16326), .B2(n16555), .C1(n16327), .C2(n16549), .A(
        n15765), .ZN(n15762) );
  AOI22_X1 U13296 ( .A1(n16545), .A2(n12436), .B1(n16537), .B2(n12308), .ZN(
        n15765) );
  OAI221_X1 U13297 ( .B1(n16321), .B2(n16555), .C1(n16322), .C2(n16549), .A(
        n15747), .ZN(n15744) );
  AOI22_X1 U13298 ( .A1(n16545), .A2(n12435), .B1(n16537), .B2(n12307), .ZN(
        n15747) );
  OAI221_X1 U13299 ( .B1(n16316), .B2(n16555), .C1(n16317), .C2(n16549), .A(
        n15729), .ZN(n15726) );
  AOI22_X1 U13300 ( .A1(n16545), .A2(n12434), .B1(n16537), .B2(n12306), .ZN(
        n15729) );
  OAI221_X1 U13301 ( .B1(n16311), .B2(n16555), .C1(n16312), .C2(n16549), .A(
        n15711), .ZN(n15708) );
  AOI22_X1 U13302 ( .A1(n16545), .A2(n12433), .B1(n16537), .B2(n12305), .ZN(
        n15711) );
  OAI221_X1 U13303 ( .B1(n16306), .B2(n16555), .C1(n16307), .C2(n16549), .A(
        n15693), .ZN(n15690) );
  AOI22_X1 U13304 ( .A1(n16545), .A2(n12432), .B1(n16537), .B2(n12304), .ZN(
        n15693) );
  OAI221_X1 U13305 ( .B1(n16301), .B2(n16555), .C1(n16302), .C2(n16549), .A(
        n15675), .ZN(n15672) );
  AOI22_X1 U13306 ( .A1(n16545), .A2(n12431), .B1(n16537), .B2(n12303), .ZN(
        n15675) );
  OAI221_X1 U13307 ( .B1(n16296), .B2(n16555), .C1(n16297), .C2(n16549), .A(
        n15657), .ZN(n15654) );
  AOI22_X1 U13308 ( .A1(n16545), .A2(n12430), .B1(n16537), .B2(n12302), .ZN(
        n15657) );
  OAI221_X1 U13309 ( .B1(n16291), .B2(n16556), .C1(n16292), .C2(n16550), .A(
        n15639), .ZN(n15636) );
  AOI22_X1 U13310 ( .A1(n16545), .A2(n12429), .B1(n16538), .B2(n12301), .ZN(
        n15639) );
  OAI221_X1 U13311 ( .B1(n16286), .B2(n16556), .C1(n16287), .C2(n16550), .A(
        n15621), .ZN(n15618) );
  AOI22_X1 U13312 ( .A1(n16545), .A2(n12428), .B1(n16538), .B2(n12300), .ZN(
        n15621) );
  OAI221_X1 U13313 ( .B1(n16281), .B2(n16556), .C1(n16282), .C2(n16550), .A(
        n15603), .ZN(n15600) );
  AOI22_X1 U13314 ( .A1(n16545), .A2(n12427), .B1(n16538), .B2(n12299), .ZN(
        n15603) );
  OAI221_X1 U13315 ( .B1(n16276), .B2(n16556), .C1(n16277), .C2(n16550), .A(
        n15585), .ZN(n15582) );
  AOI22_X1 U13316 ( .A1(n16545), .A2(n12426), .B1(n16538), .B2(n12298), .ZN(
        n15585) );
  OAI221_X1 U13317 ( .B1(n16271), .B2(n16556), .C1(n16272), .C2(n16550), .A(
        n15567), .ZN(n15564) );
  AOI22_X1 U13318 ( .A1(n16544), .A2(n12425), .B1(n16538), .B2(n12297), .ZN(
        n15567) );
  OAI221_X1 U13319 ( .B1(n16266), .B2(n16556), .C1(n16267), .C2(n16550), .A(
        n15549), .ZN(n15546) );
  AOI22_X1 U13320 ( .A1(n16544), .A2(n12424), .B1(n16538), .B2(n12296), .ZN(
        n15549) );
  OAI221_X1 U13321 ( .B1(n16261), .B2(n16556), .C1(n16262), .C2(n16550), .A(
        n15531), .ZN(n15528) );
  AOI22_X1 U13322 ( .A1(n16544), .A2(n12423), .B1(n16538), .B2(n12295), .ZN(
        n15531) );
  OAI221_X1 U13323 ( .B1(n16256), .B2(n16556), .C1(n16257), .C2(n16550), .A(
        n15513), .ZN(n15510) );
  AOI22_X1 U13324 ( .A1(n16544), .A2(n12422), .B1(n16538), .B2(n12294), .ZN(
        n15513) );
  OAI221_X1 U13325 ( .B1(n16251), .B2(n16556), .C1(n16252), .C2(n16550), .A(
        n15495), .ZN(n15492) );
  AOI22_X1 U13326 ( .A1(n16544), .A2(n12421), .B1(n16538), .B2(n12293), .ZN(
        n15495) );
  OAI221_X1 U13327 ( .B1(n16246), .B2(n16556), .C1(n16247), .C2(n16550), .A(
        n15477), .ZN(n15474) );
  AOI22_X1 U13328 ( .A1(n16544), .A2(n12420), .B1(n16538), .B2(n12292), .ZN(
        n15477) );
  OAI221_X1 U13329 ( .B1(n16241), .B2(n16556), .C1(n16242), .C2(n16550), .A(
        n15459), .ZN(n15456) );
  AOI22_X1 U13330 ( .A1(n16544), .A2(n12419), .B1(n16538), .B2(n12291), .ZN(
        n15459) );
  OAI221_X1 U13331 ( .B1(n16236), .B2(n16556), .C1(n16237), .C2(n16550), .A(
        n15441), .ZN(n15438) );
  AOI22_X1 U13332 ( .A1(n16544), .A2(n12418), .B1(n16538), .B2(n12290), .ZN(
        n15441) );
  OAI221_X1 U13333 ( .B1(n16231), .B2(n16557), .C1(n16232), .C2(n16551), .A(
        n15423), .ZN(n15420) );
  AOI22_X1 U13334 ( .A1(n16544), .A2(n12417), .B1(n16539), .B2(n12289), .ZN(
        n15423) );
  OAI221_X1 U13335 ( .B1(n16226), .B2(n16557), .C1(n16227), .C2(n16551), .A(
        n15405), .ZN(n15402) );
  AOI22_X1 U13336 ( .A1(n16544), .A2(n12416), .B1(n16539), .B2(n12288), .ZN(
        n15405) );
  OAI221_X1 U13337 ( .B1(n16221), .B2(n16557), .C1(n16222), .C2(n16551), .A(
        n15387), .ZN(n15384) );
  AOI22_X1 U13338 ( .A1(n16544), .A2(n12415), .B1(n16539), .B2(n12287), .ZN(
        n15387) );
  OAI221_X1 U13339 ( .B1(n16216), .B2(n16557), .C1(n16217), .C2(n16551), .A(
        n15369), .ZN(n15366) );
  AOI22_X1 U13340 ( .A1(n16544), .A2(n12414), .B1(n16539), .B2(n12286), .ZN(
        n15369) );
  OAI221_X1 U13341 ( .B1(n16211), .B2(n16557), .C1(n16212), .C2(n16551), .A(
        n15351), .ZN(n15348) );
  AOI22_X1 U13342 ( .A1(n16543), .A2(n12413), .B1(n16539), .B2(n12285), .ZN(
        n15351) );
  OAI221_X1 U13343 ( .B1(n16206), .B2(n16557), .C1(n16207), .C2(n16551), .A(
        n15333), .ZN(n15330) );
  AOI22_X1 U13344 ( .A1(n16543), .A2(n12412), .B1(n16539), .B2(n12284), .ZN(
        n15333) );
  OAI221_X1 U13345 ( .B1(n16201), .B2(n16557), .C1(n16202), .C2(n16551), .A(
        n15315), .ZN(n15312) );
  AOI22_X1 U13346 ( .A1(n16543), .A2(n12411), .B1(n16539), .B2(n12283), .ZN(
        n15315) );
  OAI221_X1 U13347 ( .B1(n16196), .B2(n16557), .C1(n16197), .C2(n16551), .A(
        n15297), .ZN(n15294) );
  AOI22_X1 U13348 ( .A1(n16543), .A2(n12410), .B1(n16539), .B2(n12282), .ZN(
        n15297) );
  OAI221_X1 U13349 ( .B1(n16191), .B2(n16557), .C1(n16192), .C2(n16551), .A(
        n15279), .ZN(n15276) );
  AOI22_X1 U13350 ( .A1(n16543), .A2(n12409), .B1(n16539), .B2(n12281), .ZN(
        n15279) );
  OAI221_X1 U13351 ( .B1(n16186), .B2(n16557), .C1(n16187), .C2(n16551), .A(
        n15261), .ZN(n15258) );
  AOI22_X1 U13352 ( .A1(n16543), .A2(n12408), .B1(n16539), .B2(n12280), .ZN(
        n15261) );
  OAI221_X1 U13353 ( .B1(n16181), .B2(n16557), .C1(n16182), .C2(n16551), .A(
        n15243), .ZN(n15240) );
  AOI22_X1 U13354 ( .A1(n16543), .A2(n12407), .B1(n16539), .B2(n12279), .ZN(
        n15243) );
  OAI221_X1 U13355 ( .B1(n16176), .B2(n16557), .C1(n16177), .C2(n16551), .A(
        n15225), .ZN(n15222) );
  AOI22_X1 U13356 ( .A1(n16543), .A2(n12406), .B1(n16539), .B2(n12278), .ZN(
        n15225) );
  OAI221_X1 U13357 ( .B1(n16171), .B2(n16558), .C1(n16172), .C2(n16552), .A(
        n15207), .ZN(n15204) );
  AOI22_X1 U13358 ( .A1(n16543), .A2(n12405), .B1(n16540), .B2(n12277), .ZN(
        n15207) );
  OAI221_X1 U13359 ( .B1(n16166), .B2(n16558), .C1(n16167), .C2(n16552), .A(
        n15189), .ZN(n15186) );
  AOI22_X1 U13360 ( .A1(n16543), .A2(n12404), .B1(n16540), .B2(n12276), .ZN(
        n15189) );
  OAI221_X1 U13361 ( .B1(n16161), .B2(n16558), .C1(n16162), .C2(n16552), .A(
        n15171), .ZN(n15168) );
  AOI22_X1 U13362 ( .A1(n16543), .A2(n12403), .B1(n16540), .B2(n12275), .ZN(
        n15171) );
  OAI221_X1 U13363 ( .B1(n16156), .B2(n16558), .C1(n16157), .C2(n16552), .A(
        n15153), .ZN(n15150) );
  AOI22_X1 U13364 ( .A1(n16543), .A2(n12402), .B1(n16540), .B2(n12274), .ZN(
        n15153) );
  OAI221_X1 U13365 ( .B1(n16151), .B2(n16558), .C1(n16152), .C2(n16552), .A(
        n15135), .ZN(n15132) );
  AOI22_X1 U13366 ( .A1(n16542), .A2(n12401), .B1(n16540), .B2(n12273), .ZN(
        n15135) );
  OAI221_X1 U13367 ( .B1(n16146), .B2(n16558), .C1(n16147), .C2(n16552), .A(
        n15117), .ZN(n15114) );
  AOI22_X1 U13368 ( .A1(n16542), .A2(n12400), .B1(n16540), .B2(n12272), .ZN(
        n15117) );
  OAI221_X1 U13369 ( .B1(n16141), .B2(n16558), .C1(n16142), .C2(n16552), .A(
        n15099), .ZN(n15096) );
  AOI22_X1 U13370 ( .A1(n16542), .A2(n12399), .B1(n16540), .B2(n12271), .ZN(
        n15099) );
  OAI221_X1 U13371 ( .B1(n16136), .B2(n16558), .C1(n16137), .C2(n16552), .A(
        n15081), .ZN(n15078) );
  AOI22_X1 U13372 ( .A1(n16542), .A2(n12398), .B1(n16540), .B2(n12270), .ZN(
        n15081) );
  OAI221_X1 U13373 ( .B1(n16131), .B2(n16558), .C1(n16132), .C2(n16552), .A(
        n15063), .ZN(n15060) );
  AOI22_X1 U13374 ( .A1(n16542), .A2(n12397), .B1(n16540), .B2(n12269), .ZN(
        n15063) );
  OAI221_X1 U13375 ( .B1(n16126), .B2(n16558), .C1(n16127), .C2(n16552), .A(
        n15045), .ZN(n15042) );
  AOI22_X1 U13376 ( .A1(n16542), .A2(n12396), .B1(n16540), .B2(n12268), .ZN(
        n15045) );
  OAI221_X1 U13377 ( .B1(n16121), .B2(n16558), .C1(n16122), .C2(n16552), .A(
        n15027), .ZN(n15024) );
  AOI22_X1 U13378 ( .A1(n16542), .A2(n12395), .B1(n16540), .B2(n12267), .ZN(
        n15027) );
  OAI221_X1 U13379 ( .B1(n16116), .B2(n16558), .C1(n16117), .C2(n16552), .A(
        n15009), .ZN(n15006) );
  AOI22_X1 U13380 ( .A1(n16542), .A2(n12394), .B1(n16540), .B2(n12266), .ZN(
        n15009) );
  OAI221_X1 U13381 ( .B1(n840), .B2(n16660), .C1(n12713), .C2(n16654), .A(
        n14983), .ZN(n14980) );
  AOI22_X1 U13382 ( .A1(n16648), .A2(n8188), .B1(n16642), .B2(n8252), .ZN(
        n14983) );
  OAI221_X1 U13383 ( .B1(n839), .B2(n16660), .C1(n12712), .C2(n16654), .A(
        n14965), .ZN(n14962) );
  AOI22_X1 U13384 ( .A1(n16648), .A2(n8187), .B1(n16642), .B2(n8251), .ZN(
        n14965) );
  OAI221_X1 U13385 ( .B1(n838), .B2(n16660), .C1(n12711), .C2(n16654), .A(
        n14947), .ZN(n14944) );
  AOI22_X1 U13386 ( .A1(n16648), .A2(n8186), .B1(n16642), .B2(n8250), .ZN(
        n14947) );
  OAI221_X1 U13387 ( .B1(n837), .B2(n16660), .C1(n12710), .C2(n16654), .A(
        n14901), .ZN(n14892) );
  AOI22_X1 U13388 ( .A1(n16648), .A2(n8185), .B1(n16642), .B2(n8249), .ZN(
        n14901) );
  OAI221_X1 U13389 ( .B1(n840), .B2(n16865), .C1(n12713), .C2(n16859), .A(
        n13775), .ZN(n13772) );
  AOI22_X1 U13390 ( .A1(n16853), .A2(n8188), .B1(n16847), .B2(n8252), .ZN(
        n13775) );
  OAI221_X1 U13391 ( .B1(n839), .B2(n16865), .C1(n12712), .C2(n16859), .A(
        n13757), .ZN(n13754) );
  AOI22_X1 U13392 ( .A1(n16853), .A2(n8187), .B1(n16847), .B2(n8251), .ZN(
        n13757) );
  OAI221_X1 U13393 ( .B1(n838), .B2(n16865), .C1(n12711), .C2(n16859), .A(
        n13739), .ZN(n13736) );
  AOI22_X1 U13394 ( .A1(n16853), .A2(n8186), .B1(n16847), .B2(n8250), .ZN(
        n13739) );
  OAI221_X1 U13395 ( .B1(n837), .B2(n16865), .C1(n12710), .C2(n16859), .A(
        n13693), .ZN(n13684) );
  AOI22_X1 U13396 ( .A1(n16853), .A2(n8185), .B1(n16847), .B2(n8249), .ZN(
        n13693) );
  OAI221_X1 U13397 ( .B1(n900), .B2(n16655), .C1(n12773), .C2(n16649), .A(
        n16071), .ZN(n16060) );
  AOI22_X1 U13398 ( .A1(n16643), .A2(n8248), .B1(n16637), .B2(n8312), .ZN(
        n16071) );
  OAI221_X1 U13399 ( .B1(n899), .B2(n16655), .C1(n12772), .C2(n16649), .A(
        n16045), .ZN(n16042) );
  AOI22_X1 U13400 ( .A1(n16643), .A2(n8247), .B1(n16637), .B2(n8311), .ZN(
        n16045) );
  OAI221_X1 U13401 ( .B1(n16406), .B2(n16554), .C1(n16407), .C2(n16548), .A(
        n16053), .ZN(n16050) );
  AOI22_X1 U13402 ( .A1(n16547), .A2(n12452), .B1(n16536), .B2(n12324), .ZN(
        n16053) );
  OAI221_X1 U13403 ( .B1(n898), .B2(n16655), .C1(n12771), .C2(n16649), .A(
        n16027), .ZN(n16024) );
  AOI22_X1 U13404 ( .A1(n16643), .A2(n8246), .B1(n16637), .B2(n8310), .ZN(
        n16027) );
  OAI221_X1 U13405 ( .B1(n16401), .B2(n16554), .C1(n16402), .C2(n16548), .A(
        n16035), .ZN(n16032) );
  AOI22_X1 U13406 ( .A1(n16547), .A2(n12451), .B1(n16536), .B2(n12323), .ZN(
        n16035) );
  OAI221_X1 U13407 ( .B1(n897), .B2(n16655), .C1(n12770), .C2(n16649), .A(
        n16009), .ZN(n16006) );
  AOI22_X1 U13408 ( .A1(n16643), .A2(n8245), .B1(n16637), .B2(n8309), .ZN(
        n16009) );
  OAI221_X1 U13409 ( .B1(n16396), .B2(n16554), .C1(n16397), .C2(n16548), .A(
        n16017), .ZN(n16014) );
  AOI22_X1 U13410 ( .A1(n16547), .A2(n12450), .B1(n16536), .B2(n12322), .ZN(
        n16017) );
  OAI221_X1 U13411 ( .B1(n896), .B2(n16655), .C1(n12769), .C2(n16649), .A(
        n15991), .ZN(n15988) );
  AOI22_X1 U13412 ( .A1(n16643), .A2(n8244), .B1(n16637), .B2(n8308), .ZN(
        n15991) );
  OAI221_X1 U13413 ( .B1(n16391), .B2(n16554), .C1(n16392), .C2(n16548), .A(
        n15999), .ZN(n15996) );
  AOI22_X1 U13414 ( .A1(n16546), .A2(n12449), .B1(n16536), .B2(n12321), .ZN(
        n15999) );
  OAI221_X1 U13415 ( .B1(n895), .B2(n16655), .C1(n12768), .C2(n16649), .A(
        n15973), .ZN(n15970) );
  AOI22_X1 U13416 ( .A1(n16643), .A2(n8243), .B1(n16637), .B2(n8307), .ZN(
        n15973) );
  OAI221_X1 U13417 ( .B1(n16386), .B2(n16554), .C1(n16387), .C2(n16548), .A(
        n15981), .ZN(n15978) );
  AOI22_X1 U13418 ( .A1(n16546), .A2(n12448), .B1(n16536), .B2(n12320), .ZN(
        n15981) );
  OAI221_X1 U13419 ( .B1(n894), .B2(n16655), .C1(n12767), .C2(n16649), .A(
        n15955), .ZN(n15952) );
  AOI22_X1 U13420 ( .A1(n16643), .A2(n8242), .B1(n16637), .B2(n8306), .ZN(
        n15955) );
  OAI221_X1 U13421 ( .B1(n16381), .B2(n16554), .C1(n16382), .C2(n16548), .A(
        n15963), .ZN(n15960) );
  AOI22_X1 U13422 ( .A1(n16546), .A2(n12447), .B1(n16536), .B2(n12319), .ZN(
        n15963) );
  OAI221_X1 U13423 ( .B1(n893), .B2(n16655), .C1(n12766), .C2(n16649), .A(
        n15937), .ZN(n15934) );
  AOI22_X1 U13424 ( .A1(n16643), .A2(n8241), .B1(n16637), .B2(n8305), .ZN(
        n15937) );
  OAI221_X1 U13425 ( .B1(n16376), .B2(n16554), .C1(n16377), .C2(n16548), .A(
        n15945), .ZN(n15942) );
  AOI22_X1 U13426 ( .A1(n16546), .A2(n12446), .B1(n16536), .B2(n12318), .ZN(
        n15945) );
  OAI221_X1 U13427 ( .B1(n892), .B2(n16655), .C1(n12765), .C2(n16649), .A(
        n15919), .ZN(n15916) );
  AOI22_X1 U13428 ( .A1(n16643), .A2(n8240), .B1(n16637), .B2(n8304), .ZN(
        n15919) );
  OAI221_X1 U13429 ( .B1(n16371), .B2(n16554), .C1(n16372), .C2(n16548), .A(
        n15927), .ZN(n15924) );
  AOI22_X1 U13430 ( .A1(n16546), .A2(n12445), .B1(n16536), .B2(n12317), .ZN(
        n15927) );
  OAI221_X1 U13431 ( .B1(n891), .B2(n16655), .C1(n12764), .C2(n16649), .A(
        n15901), .ZN(n15898) );
  AOI22_X1 U13432 ( .A1(n16643), .A2(n8239), .B1(n16637), .B2(n8303), .ZN(
        n15901) );
  OAI221_X1 U13433 ( .B1(n16366), .B2(n16554), .C1(n16367), .C2(n16548), .A(
        n15909), .ZN(n15906) );
  AOI22_X1 U13434 ( .A1(n16546), .A2(n12444), .B1(n16536), .B2(n12316), .ZN(
        n15909) );
  OAI221_X1 U13435 ( .B1(n890), .B2(n16655), .C1(n12763), .C2(n16649), .A(
        n15883), .ZN(n15880) );
  AOI22_X1 U13436 ( .A1(n16643), .A2(n8238), .B1(n16637), .B2(n8302), .ZN(
        n15883) );
  OAI221_X1 U13437 ( .B1(n16361), .B2(n16554), .C1(n16362), .C2(n16548), .A(
        n15891), .ZN(n15888) );
  AOI22_X1 U13438 ( .A1(n16546), .A2(n12443), .B1(n16536), .B2(n12315), .ZN(
        n15891) );
  OAI221_X1 U13439 ( .B1(n889), .B2(n16655), .C1(n12762), .C2(n16649), .A(
        n15865), .ZN(n15862) );
  AOI22_X1 U13440 ( .A1(n16643), .A2(n8237), .B1(n16637), .B2(n8301), .ZN(
        n15865) );
  OAI221_X1 U13441 ( .B1(n16356), .B2(n16554), .C1(n16357), .C2(n16548), .A(
        n15873), .ZN(n15870) );
  AOI22_X1 U13442 ( .A1(n16546), .A2(n12442), .B1(n16536), .B2(n12314), .ZN(
        n15873) );
  OAI221_X1 U13443 ( .B1(n888), .B2(n16656), .C1(n12761), .C2(n16650), .A(
        n15847), .ZN(n15844) );
  AOI22_X1 U13444 ( .A1(n16644), .A2(n8236), .B1(n16638), .B2(n8300), .ZN(
        n15847) );
  OAI221_X1 U13445 ( .B1(n887), .B2(n16656), .C1(n12760), .C2(n16650), .A(
        n15829), .ZN(n15826) );
  AOI22_X1 U13446 ( .A1(n16644), .A2(n8235), .B1(n16638), .B2(n8299), .ZN(
        n15829) );
  OAI221_X1 U13447 ( .B1(n886), .B2(n16656), .C1(n12759), .C2(n16650), .A(
        n15811), .ZN(n15808) );
  AOI22_X1 U13448 ( .A1(n16644), .A2(n8234), .B1(n16638), .B2(n8298), .ZN(
        n15811) );
  OAI221_X1 U13449 ( .B1(n885), .B2(n16656), .C1(n12758), .C2(n16650), .A(
        n15793), .ZN(n15790) );
  AOI22_X1 U13450 ( .A1(n16644), .A2(n8233), .B1(n16638), .B2(n8297), .ZN(
        n15793) );
  OAI221_X1 U13451 ( .B1(n884), .B2(n16656), .C1(n12757), .C2(n16650), .A(
        n15775), .ZN(n15772) );
  AOI22_X1 U13452 ( .A1(n16644), .A2(n8232), .B1(n16638), .B2(n8296), .ZN(
        n15775) );
  OAI221_X1 U13453 ( .B1(n883), .B2(n16656), .C1(n12756), .C2(n16650), .A(
        n15757), .ZN(n15754) );
  AOI22_X1 U13454 ( .A1(n16644), .A2(n8231), .B1(n16638), .B2(n8295), .ZN(
        n15757) );
  OAI221_X1 U13455 ( .B1(n882), .B2(n16656), .C1(n12755), .C2(n16650), .A(
        n15739), .ZN(n15736) );
  AOI22_X1 U13456 ( .A1(n16644), .A2(n8230), .B1(n16638), .B2(n8294), .ZN(
        n15739) );
  OAI221_X1 U13457 ( .B1(n881), .B2(n16656), .C1(n12754), .C2(n16650), .A(
        n15721), .ZN(n15718) );
  AOI22_X1 U13458 ( .A1(n16644), .A2(n8229), .B1(n16638), .B2(n8293), .ZN(
        n15721) );
  OAI221_X1 U13459 ( .B1(n880), .B2(n16656), .C1(n12753), .C2(n16650), .A(
        n15703), .ZN(n15700) );
  AOI22_X1 U13460 ( .A1(n16644), .A2(n8228), .B1(n16638), .B2(n8292), .ZN(
        n15703) );
  OAI221_X1 U13461 ( .B1(n879), .B2(n16656), .C1(n12752), .C2(n16650), .A(
        n15685), .ZN(n15682) );
  AOI22_X1 U13462 ( .A1(n16644), .A2(n8227), .B1(n16638), .B2(n8291), .ZN(
        n15685) );
  OAI221_X1 U13463 ( .B1(n878), .B2(n16656), .C1(n12751), .C2(n16650), .A(
        n15667), .ZN(n15664) );
  AOI22_X1 U13464 ( .A1(n16644), .A2(n8226), .B1(n16638), .B2(n8290), .ZN(
        n15667) );
  OAI221_X1 U13465 ( .B1(n877), .B2(n16656), .C1(n12750), .C2(n16650), .A(
        n15649), .ZN(n15646) );
  AOI22_X1 U13466 ( .A1(n16644), .A2(n8225), .B1(n16638), .B2(n8289), .ZN(
        n15649) );
  OAI221_X1 U13467 ( .B1(n876), .B2(n16657), .C1(n12749), .C2(n16651), .A(
        n15631), .ZN(n15628) );
  AOI22_X1 U13468 ( .A1(n16645), .A2(n8224), .B1(n16639), .B2(n8288), .ZN(
        n15631) );
  OAI221_X1 U13469 ( .B1(n875), .B2(n16657), .C1(n12748), .C2(n16651), .A(
        n15613), .ZN(n15610) );
  AOI22_X1 U13470 ( .A1(n16645), .A2(n8223), .B1(n16639), .B2(n8287), .ZN(
        n15613) );
  OAI221_X1 U13471 ( .B1(n874), .B2(n16657), .C1(n12747), .C2(n16651), .A(
        n15595), .ZN(n15592) );
  AOI22_X1 U13472 ( .A1(n16645), .A2(n8222), .B1(n16639), .B2(n8286), .ZN(
        n15595) );
  OAI221_X1 U13473 ( .B1(n873), .B2(n16657), .C1(n12746), .C2(n16651), .A(
        n15577), .ZN(n15574) );
  AOI22_X1 U13474 ( .A1(n16645), .A2(n8221), .B1(n16639), .B2(n8285), .ZN(
        n15577) );
  OAI221_X1 U13475 ( .B1(n872), .B2(n16657), .C1(n12745), .C2(n16651), .A(
        n15559), .ZN(n15556) );
  AOI22_X1 U13476 ( .A1(n16645), .A2(n8220), .B1(n16639), .B2(n8284), .ZN(
        n15559) );
  OAI221_X1 U13477 ( .B1(n871), .B2(n16657), .C1(n12744), .C2(n16651), .A(
        n15541), .ZN(n15538) );
  AOI22_X1 U13478 ( .A1(n16645), .A2(n8219), .B1(n16639), .B2(n8283), .ZN(
        n15541) );
  OAI221_X1 U13479 ( .B1(n870), .B2(n16657), .C1(n12743), .C2(n16651), .A(
        n15523), .ZN(n15520) );
  AOI22_X1 U13480 ( .A1(n16645), .A2(n8218), .B1(n16639), .B2(n8282), .ZN(
        n15523) );
  OAI221_X1 U13481 ( .B1(n869), .B2(n16657), .C1(n12742), .C2(n16651), .A(
        n15505), .ZN(n15502) );
  AOI22_X1 U13482 ( .A1(n16645), .A2(n8217), .B1(n16639), .B2(n8281), .ZN(
        n15505) );
  OAI221_X1 U13483 ( .B1(n868), .B2(n16657), .C1(n12741), .C2(n16651), .A(
        n15487), .ZN(n15484) );
  AOI22_X1 U13484 ( .A1(n16645), .A2(n8216), .B1(n16639), .B2(n8280), .ZN(
        n15487) );
  OAI221_X1 U13485 ( .B1(n867), .B2(n16657), .C1(n12740), .C2(n16651), .A(
        n15469), .ZN(n15466) );
  AOI22_X1 U13486 ( .A1(n16645), .A2(n8215), .B1(n16639), .B2(n8279), .ZN(
        n15469) );
  OAI221_X1 U13487 ( .B1(n866), .B2(n16657), .C1(n12739), .C2(n16651), .A(
        n15451), .ZN(n15448) );
  AOI22_X1 U13488 ( .A1(n16645), .A2(n8214), .B1(n16639), .B2(n8278), .ZN(
        n15451) );
  OAI221_X1 U13489 ( .B1(n865), .B2(n16657), .C1(n12738), .C2(n16651), .A(
        n15433), .ZN(n15430) );
  AOI22_X1 U13490 ( .A1(n16645), .A2(n8213), .B1(n16639), .B2(n8277), .ZN(
        n15433) );
  OAI221_X1 U13491 ( .B1(n864), .B2(n16658), .C1(n12737), .C2(n16652), .A(
        n15415), .ZN(n15412) );
  AOI22_X1 U13492 ( .A1(n16646), .A2(n8212), .B1(n16640), .B2(n8276), .ZN(
        n15415) );
  OAI221_X1 U13493 ( .B1(n863), .B2(n16658), .C1(n12736), .C2(n16652), .A(
        n15397), .ZN(n15394) );
  AOI22_X1 U13494 ( .A1(n16646), .A2(n8211), .B1(n16640), .B2(n8275), .ZN(
        n15397) );
  OAI221_X1 U13495 ( .B1(n862), .B2(n16658), .C1(n12735), .C2(n16652), .A(
        n15379), .ZN(n15376) );
  AOI22_X1 U13496 ( .A1(n16646), .A2(n8210), .B1(n16640), .B2(n8274), .ZN(
        n15379) );
  OAI221_X1 U13497 ( .B1(n861), .B2(n16658), .C1(n12734), .C2(n16652), .A(
        n15361), .ZN(n15358) );
  AOI22_X1 U13498 ( .A1(n16646), .A2(n8209), .B1(n16640), .B2(n8273), .ZN(
        n15361) );
  OAI221_X1 U13499 ( .B1(n860), .B2(n16658), .C1(n12733), .C2(n16652), .A(
        n15343), .ZN(n15340) );
  AOI22_X1 U13500 ( .A1(n16646), .A2(n8208), .B1(n16640), .B2(n8272), .ZN(
        n15343) );
  OAI221_X1 U13501 ( .B1(n859), .B2(n16658), .C1(n12732), .C2(n16652), .A(
        n15325), .ZN(n15322) );
  AOI22_X1 U13502 ( .A1(n16646), .A2(n8207), .B1(n16640), .B2(n8271), .ZN(
        n15325) );
  OAI221_X1 U13503 ( .B1(n858), .B2(n16658), .C1(n12731), .C2(n16652), .A(
        n15307), .ZN(n15304) );
  AOI22_X1 U13504 ( .A1(n16646), .A2(n8206), .B1(n16640), .B2(n8270), .ZN(
        n15307) );
  OAI221_X1 U13505 ( .B1(n857), .B2(n16658), .C1(n12730), .C2(n16652), .A(
        n15289), .ZN(n15286) );
  AOI22_X1 U13506 ( .A1(n16646), .A2(n8205), .B1(n16640), .B2(n8269), .ZN(
        n15289) );
  OAI221_X1 U13507 ( .B1(n856), .B2(n16658), .C1(n12729), .C2(n16652), .A(
        n15271), .ZN(n15268) );
  AOI22_X1 U13508 ( .A1(n16646), .A2(n8204), .B1(n16640), .B2(n8268), .ZN(
        n15271) );
  OAI221_X1 U13509 ( .B1(n855), .B2(n16658), .C1(n12728), .C2(n16652), .A(
        n15253), .ZN(n15250) );
  AOI22_X1 U13510 ( .A1(n16646), .A2(n8203), .B1(n16640), .B2(n8267), .ZN(
        n15253) );
  OAI221_X1 U13511 ( .B1(n854), .B2(n16658), .C1(n12727), .C2(n16652), .A(
        n15235), .ZN(n15232) );
  AOI22_X1 U13512 ( .A1(n16646), .A2(n8202), .B1(n16640), .B2(n8266), .ZN(
        n15235) );
  OAI221_X1 U13513 ( .B1(n853), .B2(n16658), .C1(n12726), .C2(n16652), .A(
        n15217), .ZN(n15214) );
  AOI22_X1 U13514 ( .A1(n16646), .A2(n8201), .B1(n16640), .B2(n8265), .ZN(
        n15217) );
  OAI221_X1 U13515 ( .B1(n852), .B2(n16659), .C1(n12725), .C2(n16653), .A(
        n15199), .ZN(n15196) );
  AOI22_X1 U13516 ( .A1(n16647), .A2(n8200), .B1(n16641), .B2(n8264), .ZN(
        n15199) );
  OAI221_X1 U13517 ( .B1(n851), .B2(n16659), .C1(n12724), .C2(n16653), .A(
        n15181), .ZN(n15178) );
  AOI22_X1 U13518 ( .A1(n16647), .A2(n8199), .B1(n16641), .B2(n8263), .ZN(
        n15181) );
  OAI221_X1 U13519 ( .B1(n850), .B2(n16659), .C1(n12723), .C2(n16653), .A(
        n15163), .ZN(n15160) );
  AOI22_X1 U13520 ( .A1(n16647), .A2(n8198), .B1(n16641), .B2(n8262), .ZN(
        n15163) );
  OAI221_X1 U13521 ( .B1(n849), .B2(n16659), .C1(n12722), .C2(n16653), .A(
        n15145), .ZN(n15142) );
  AOI22_X1 U13522 ( .A1(n16647), .A2(n8197), .B1(n16641), .B2(n8261), .ZN(
        n15145) );
  OAI221_X1 U13523 ( .B1(n848), .B2(n16659), .C1(n12721), .C2(n16653), .A(
        n15127), .ZN(n15124) );
  AOI22_X1 U13524 ( .A1(n16647), .A2(n8196), .B1(n16641), .B2(n8260), .ZN(
        n15127) );
  OAI221_X1 U13525 ( .B1(n847), .B2(n16659), .C1(n12720), .C2(n16653), .A(
        n15109), .ZN(n15106) );
  AOI22_X1 U13526 ( .A1(n16647), .A2(n8195), .B1(n16641), .B2(n8259), .ZN(
        n15109) );
  OAI221_X1 U13527 ( .B1(n846), .B2(n16659), .C1(n12719), .C2(n16653), .A(
        n15091), .ZN(n15088) );
  AOI22_X1 U13528 ( .A1(n16647), .A2(n8194), .B1(n16641), .B2(n8258), .ZN(
        n15091) );
  OAI221_X1 U13529 ( .B1(n845), .B2(n16659), .C1(n12718), .C2(n16653), .A(
        n15073), .ZN(n15070) );
  AOI22_X1 U13530 ( .A1(n16647), .A2(n8193), .B1(n16641), .B2(n8257), .ZN(
        n15073) );
  OAI221_X1 U13531 ( .B1(n844), .B2(n16659), .C1(n12717), .C2(n16653), .A(
        n15055), .ZN(n15052) );
  AOI22_X1 U13532 ( .A1(n16647), .A2(n8192), .B1(n16641), .B2(n8256), .ZN(
        n15055) );
  OAI221_X1 U13533 ( .B1(n843), .B2(n16659), .C1(n12716), .C2(n16653), .A(
        n15037), .ZN(n15034) );
  AOI22_X1 U13534 ( .A1(n16647), .A2(n8191), .B1(n16641), .B2(n8255), .ZN(
        n15037) );
  OAI221_X1 U13535 ( .B1(n842), .B2(n16659), .C1(n12715), .C2(n16653), .A(
        n15019), .ZN(n15016) );
  AOI22_X1 U13536 ( .A1(n16647), .A2(n8190), .B1(n16641), .B2(n8254), .ZN(
        n15019) );
  OAI221_X1 U13537 ( .B1(n841), .B2(n16659), .C1(n12714), .C2(n16653), .A(
        n15001), .ZN(n14998) );
  AOI22_X1 U13538 ( .A1(n16647), .A2(n8189), .B1(n16641), .B2(n8253), .ZN(
        n15001) );
  OAI221_X1 U13539 ( .B1(n900), .B2(n16860), .C1(n12773), .C2(n16854), .A(
        n14863), .ZN(n14852) );
  AOI22_X1 U13540 ( .A1(n16848), .A2(n8248), .B1(n16842), .B2(n8312), .ZN(
        n14863) );
  OAI221_X1 U13541 ( .B1(n899), .B2(n16860), .C1(n12772), .C2(n16854), .A(
        n14837), .ZN(n14834) );
  AOI22_X1 U13542 ( .A1(n16848), .A2(n8247), .B1(n16842), .B2(n8311), .ZN(
        n14837) );
  OAI221_X1 U13543 ( .B1(n898), .B2(n16860), .C1(n12771), .C2(n16854), .A(
        n14819), .ZN(n14816) );
  AOI22_X1 U13544 ( .A1(n16848), .A2(n8246), .B1(n16842), .B2(n8310), .ZN(
        n14819) );
  OAI221_X1 U13545 ( .B1(n897), .B2(n16860), .C1(n12770), .C2(n16854), .A(
        n14801), .ZN(n14798) );
  AOI22_X1 U13546 ( .A1(n16848), .A2(n8245), .B1(n16842), .B2(n8309), .ZN(
        n14801) );
  OAI221_X1 U13547 ( .B1(n896), .B2(n16860), .C1(n12769), .C2(n16854), .A(
        n14783), .ZN(n14780) );
  AOI22_X1 U13548 ( .A1(n16848), .A2(n8244), .B1(n16842), .B2(n8308), .ZN(
        n14783) );
  OAI221_X1 U13549 ( .B1(n895), .B2(n16860), .C1(n12768), .C2(n16854), .A(
        n14765), .ZN(n14762) );
  AOI22_X1 U13550 ( .A1(n16848), .A2(n8243), .B1(n16842), .B2(n8307), .ZN(
        n14765) );
  OAI221_X1 U13551 ( .B1(n894), .B2(n16860), .C1(n12767), .C2(n16854), .A(
        n14747), .ZN(n14744) );
  AOI22_X1 U13552 ( .A1(n16848), .A2(n8242), .B1(n16842), .B2(n8306), .ZN(
        n14747) );
  OAI221_X1 U13553 ( .B1(n893), .B2(n16860), .C1(n12766), .C2(n16854), .A(
        n14729), .ZN(n14726) );
  AOI22_X1 U13554 ( .A1(n16848), .A2(n8241), .B1(n16842), .B2(n8305), .ZN(
        n14729) );
  OAI221_X1 U13555 ( .B1(n892), .B2(n16860), .C1(n12765), .C2(n16854), .A(
        n14711), .ZN(n14708) );
  AOI22_X1 U13556 ( .A1(n16848), .A2(n8240), .B1(n16842), .B2(n8304), .ZN(
        n14711) );
  OAI221_X1 U13557 ( .B1(n891), .B2(n16860), .C1(n12764), .C2(n16854), .A(
        n14693), .ZN(n14690) );
  AOI22_X1 U13558 ( .A1(n16848), .A2(n8239), .B1(n16842), .B2(n8303), .ZN(
        n14693) );
  OAI221_X1 U13559 ( .B1(n890), .B2(n16860), .C1(n12763), .C2(n16854), .A(
        n14675), .ZN(n14672) );
  AOI22_X1 U13560 ( .A1(n16848), .A2(n8238), .B1(n16842), .B2(n8302), .ZN(
        n14675) );
  OAI221_X1 U13561 ( .B1(n889), .B2(n16860), .C1(n12762), .C2(n16854), .A(
        n14657), .ZN(n14654) );
  AOI22_X1 U13562 ( .A1(n16848), .A2(n8237), .B1(n16842), .B2(n8301), .ZN(
        n14657) );
  OAI221_X1 U13563 ( .B1(n888), .B2(n16861), .C1(n12761), .C2(n16855), .A(
        n14639), .ZN(n14636) );
  AOI22_X1 U13564 ( .A1(n16849), .A2(n8236), .B1(n16843), .B2(n8300), .ZN(
        n14639) );
  OAI221_X1 U13565 ( .B1(n887), .B2(n16861), .C1(n12760), .C2(n16855), .A(
        n14621), .ZN(n14618) );
  AOI22_X1 U13566 ( .A1(n16849), .A2(n8235), .B1(n16843), .B2(n8299), .ZN(
        n14621) );
  OAI221_X1 U13567 ( .B1(n886), .B2(n16861), .C1(n12759), .C2(n16855), .A(
        n14603), .ZN(n14600) );
  AOI22_X1 U13568 ( .A1(n16849), .A2(n8234), .B1(n16843), .B2(n8298), .ZN(
        n14603) );
  OAI221_X1 U13569 ( .B1(n885), .B2(n16861), .C1(n12758), .C2(n16855), .A(
        n14585), .ZN(n14582) );
  AOI22_X1 U13570 ( .A1(n16849), .A2(n8233), .B1(n16843), .B2(n8297), .ZN(
        n14585) );
  OAI221_X1 U13571 ( .B1(n884), .B2(n16861), .C1(n12757), .C2(n16855), .A(
        n14567), .ZN(n14564) );
  AOI22_X1 U13572 ( .A1(n16849), .A2(n8232), .B1(n16843), .B2(n8296), .ZN(
        n14567) );
  OAI221_X1 U13573 ( .B1(n883), .B2(n16861), .C1(n12756), .C2(n16855), .A(
        n14549), .ZN(n14546) );
  AOI22_X1 U13574 ( .A1(n16849), .A2(n8231), .B1(n16843), .B2(n8295), .ZN(
        n14549) );
  OAI221_X1 U13575 ( .B1(n882), .B2(n16861), .C1(n12755), .C2(n16855), .A(
        n14531), .ZN(n14528) );
  AOI22_X1 U13576 ( .A1(n16849), .A2(n8230), .B1(n16843), .B2(n8294), .ZN(
        n14531) );
  OAI221_X1 U13577 ( .B1(n881), .B2(n16861), .C1(n12754), .C2(n16855), .A(
        n14513), .ZN(n14510) );
  AOI22_X1 U13578 ( .A1(n16849), .A2(n8229), .B1(n16843), .B2(n8293), .ZN(
        n14513) );
  OAI221_X1 U13579 ( .B1(n880), .B2(n16861), .C1(n12753), .C2(n16855), .A(
        n14495), .ZN(n14492) );
  AOI22_X1 U13580 ( .A1(n16849), .A2(n8228), .B1(n16843), .B2(n8292), .ZN(
        n14495) );
  OAI221_X1 U13581 ( .B1(n879), .B2(n16861), .C1(n12752), .C2(n16855), .A(
        n14477), .ZN(n14474) );
  AOI22_X1 U13582 ( .A1(n16849), .A2(n8227), .B1(n16843), .B2(n8291), .ZN(
        n14477) );
  OAI221_X1 U13583 ( .B1(n878), .B2(n16861), .C1(n12751), .C2(n16855), .A(
        n14459), .ZN(n14456) );
  AOI22_X1 U13584 ( .A1(n16849), .A2(n8226), .B1(n16843), .B2(n8290), .ZN(
        n14459) );
  OAI221_X1 U13585 ( .B1(n877), .B2(n16861), .C1(n12750), .C2(n16855), .A(
        n14441), .ZN(n14438) );
  AOI22_X1 U13586 ( .A1(n16849), .A2(n8225), .B1(n16843), .B2(n8289), .ZN(
        n14441) );
  OAI221_X1 U13587 ( .B1(n876), .B2(n16862), .C1(n12749), .C2(n16856), .A(
        n14423), .ZN(n14420) );
  AOI22_X1 U13588 ( .A1(n16850), .A2(n8224), .B1(n16844), .B2(n8288), .ZN(
        n14423) );
  OAI221_X1 U13589 ( .B1(n875), .B2(n16862), .C1(n12748), .C2(n16856), .A(
        n14405), .ZN(n14402) );
  AOI22_X1 U13590 ( .A1(n16850), .A2(n8223), .B1(n16844), .B2(n8287), .ZN(
        n14405) );
  OAI221_X1 U13591 ( .B1(n874), .B2(n16862), .C1(n12747), .C2(n16856), .A(
        n14387), .ZN(n14384) );
  AOI22_X1 U13592 ( .A1(n16850), .A2(n8222), .B1(n16844), .B2(n8286), .ZN(
        n14387) );
  OAI221_X1 U13593 ( .B1(n873), .B2(n16862), .C1(n12746), .C2(n16856), .A(
        n14369), .ZN(n14366) );
  AOI22_X1 U13594 ( .A1(n16850), .A2(n8221), .B1(n16844), .B2(n8285), .ZN(
        n14369) );
  OAI221_X1 U13595 ( .B1(n872), .B2(n16862), .C1(n12745), .C2(n16856), .A(
        n14351), .ZN(n14348) );
  AOI22_X1 U13596 ( .A1(n16850), .A2(n8220), .B1(n16844), .B2(n8284), .ZN(
        n14351) );
  OAI221_X1 U13597 ( .B1(n871), .B2(n16862), .C1(n12744), .C2(n16856), .A(
        n14333), .ZN(n14330) );
  AOI22_X1 U13598 ( .A1(n16850), .A2(n8219), .B1(n16844), .B2(n8283), .ZN(
        n14333) );
  OAI221_X1 U13599 ( .B1(n870), .B2(n16862), .C1(n12743), .C2(n16856), .A(
        n14315), .ZN(n14312) );
  AOI22_X1 U13600 ( .A1(n16850), .A2(n8218), .B1(n16844), .B2(n8282), .ZN(
        n14315) );
  OAI221_X1 U13601 ( .B1(n869), .B2(n16862), .C1(n12742), .C2(n16856), .A(
        n14297), .ZN(n14294) );
  AOI22_X1 U13602 ( .A1(n16850), .A2(n8217), .B1(n16844), .B2(n8281), .ZN(
        n14297) );
  OAI221_X1 U13603 ( .B1(n868), .B2(n16862), .C1(n12741), .C2(n16856), .A(
        n14279), .ZN(n14276) );
  AOI22_X1 U13604 ( .A1(n16850), .A2(n8216), .B1(n16844), .B2(n8280), .ZN(
        n14279) );
  OAI221_X1 U13605 ( .B1(n867), .B2(n16862), .C1(n12740), .C2(n16856), .A(
        n14261), .ZN(n14258) );
  AOI22_X1 U13606 ( .A1(n16850), .A2(n8215), .B1(n16844), .B2(n8279), .ZN(
        n14261) );
  OAI221_X1 U13607 ( .B1(n866), .B2(n16862), .C1(n12739), .C2(n16856), .A(
        n14243), .ZN(n14240) );
  AOI22_X1 U13608 ( .A1(n16850), .A2(n8214), .B1(n16844), .B2(n8278), .ZN(
        n14243) );
  OAI221_X1 U13609 ( .B1(n865), .B2(n16862), .C1(n12738), .C2(n16856), .A(
        n14225), .ZN(n14222) );
  AOI22_X1 U13610 ( .A1(n16850), .A2(n8213), .B1(n16844), .B2(n8277), .ZN(
        n14225) );
  OAI221_X1 U13611 ( .B1(n864), .B2(n16863), .C1(n12737), .C2(n16857), .A(
        n14207), .ZN(n14204) );
  AOI22_X1 U13612 ( .A1(n16851), .A2(n8212), .B1(n16845), .B2(n8276), .ZN(
        n14207) );
  OAI221_X1 U13613 ( .B1(n863), .B2(n16863), .C1(n12736), .C2(n16857), .A(
        n14189), .ZN(n14186) );
  AOI22_X1 U13614 ( .A1(n16851), .A2(n8211), .B1(n16845), .B2(n8275), .ZN(
        n14189) );
  OAI221_X1 U13615 ( .B1(n862), .B2(n16863), .C1(n12735), .C2(n16857), .A(
        n14171), .ZN(n14168) );
  AOI22_X1 U13616 ( .A1(n16851), .A2(n8210), .B1(n16845), .B2(n8274), .ZN(
        n14171) );
  OAI221_X1 U13617 ( .B1(n861), .B2(n16863), .C1(n12734), .C2(n16857), .A(
        n14153), .ZN(n14150) );
  AOI22_X1 U13618 ( .A1(n16851), .A2(n8209), .B1(n16845), .B2(n8273), .ZN(
        n14153) );
  OAI221_X1 U13619 ( .B1(n860), .B2(n16863), .C1(n12733), .C2(n16857), .A(
        n14135), .ZN(n14132) );
  AOI22_X1 U13620 ( .A1(n16851), .A2(n8208), .B1(n16845), .B2(n8272), .ZN(
        n14135) );
  OAI221_X1 U13621 ( .B1(n859), .B2(n16863), .C1(n12732), .C2(n16857), .A(
        n14117), .ZN(n14114) );
  AOI22_X1 U13622 ( .A1(n16851), .A2(n8207), .B1(n16845), .B2(n8271), .ZN(
        n14117) );
  OAI221_X1 U13623 ( .B1(n858), .B2(n16863), .C1(n12731), .C2(n16857), .A(
        n14099), .ZN(n14096) );
  AOI22_X1 U13624 ( .A1(n16851), .A2(n8206), .B1(n16845), .B2(n8270), .ZN(
        n14099) );
  OAI221_X1 U13625 ( .B1(n857), .B2(n16863), .C1(n12730), .C2(n16857), .A(
        n14081), .ZN(n14078) );
  AOI22_X1 U13626 ( .A1(n16851), .A2(n8205), .B1(n16845), .B2(n8269), .ZN(
        n14081) );
  OAI221_X1 U13627 ( .B1(n856), .B2(n16863), .C1(n12729), .C2(n16857), .A(
        n14063), .ZN(n14060) );
  AOI22_X1 U13628 ( .A1(n16851), .A2(n8204), .B1(n16845), .B2(n8268), .ZN(
        n14063) );
  OAI221_X1 U13629 ( .B1(n855), .B2(n16863), .C1(n12728), .C2(n16857), .A(
        n14045), .ZN(n14042) );
  AOI22_X1 U13630 ( .A1(n16851), .A2(n8203), .B1(n16845), .B2(n8267), .ZN(
        n14045) );
  OAI221_X1 U13631 ( .B1(n854), .B2(n16863), .C1(n12727), .C2(n16857), .A(
        n14027), .ZN(n14024) );
  AOI22_X1 U13632 ( .A1(n16851), .A2(n8202), .B1(n16845), .B2(n8266), .ZN(
        n14027) );
  OAI221_X1 U13633 ( .B1(n853), .B2(n16863), .C1(n12726), .C2(n16857), .A(
        n14009), .ZN(n14006) );
  AOI22_X1 U13634 ( .A1(n16851), .A2(n8201), .B1(n16845), .B2(n8265), .ZN(
        n14009) );
  OAI221_X1 U13635 ( .B1(n852), .B2(n16864), .C1(n12725), .C2(n16858), .A(
        n13991), .ZN(n13988) );
  AOI22_X1 U13636 ( .A1(n16852), .A2(n8200), .B1(n16846), .B2(n8264), .ZN(
        n13991) );
  OAI221_X1 U13637 ( .B1(n851), .B2(n16864), .C1(n12724), .C2(n16858), .A(
        n13973), .ZN(n13970) );
  AOI22_X1 U13638 ( .A1(n16852), .A2(n8199), .B1(n16846), .B2(n8263), .ZN(
        n13973) );
  OAI221_X1 U13639 ( .B1(n850), .B2(n16864), .C1(n12723), .C2(n16858), .A(
        n13955), .ZN(n13952) );
  AOI22_X1 U13640 ( .A1(n16852), .A2(n8198), .B1(n16846), .B2(n8262), .ZN(
        n13955) );
  OAI221_X1 U13641 ( .B1(n849), .B2(n16864), .C1(n12722), .C2(n16858), .A(
        n13937), .ZN(n13934) );
  AOI22_X1 U13642 ( .A1(n16852), .A2(n8197), .B1(n16846), .B2(n8261), .ZN(
        n13937) );
  OAI221_X1 U13643 ( .B1(n848), .B2(n16864), .C1(n12721), .C2(n16858), .A(
        n13919), .ZN(n13916) );
  AOI22_X1 U13644 ( .A1(n16852), .A2(n8196), .B1(n16846), .B2(n8260), .ZN(
        n13919) );
  OAI221_X1 U13645 ( .B1(n847), .B2(n16864), .C1(n12720), .C2(n16858), .A(
        n13901), .ZN(n13898) );
  AOI22_X1 U13646 ( .A1(n16852), .A2(n8195), .B1(n16846), .B2(n8259), .ZN(
        n13901) );
  OAI221_X1 U13647 ( .B1(n846), .B2(n16864), .C1(n12719), .C2(n16858), .A(
        n13883), .ZN(n13880) );
  AOI22_X1 U13648 ( .A1(n16852), .A2(n8194), .B1(n16846), .B2(n8258), .ZN(
        n13883) );
  OAI221_X1 U13649 ( .B1(n845), .B2(n16864), .C1(n12718), .C2(n16858), .A(
        n13865), .ZN(n13862) );
  AOI22_X1 U13650 ( .A1(n16852), .A2(n8193), .B1(n16846), .B2(n8257), .ZN(
        n13865) );
  OAI221_X1 U13651 ( .B1(n844), .B2(n16864), .C1(n12717), .C2(n16858), .A(
        n13847), .ZN(n13844) );
  AOI22_X1 U13652 ( .A1(n16852), .A2(n8192), .B1(n16846), .B2(n8256), .ZN(
        n13847) );
  OAI221_X1 U13653 ( .B1(n843), .B2(n16864), .C1(n12716), .C2(n16858), .A(
        n13829), .ZN(n13826) );
  AOI22_X1 U13654 ( .A1(n16852), .A2(n8191), .B1(n16846), .B2(n8255), .ZN(
        n13829) );
  OAI221_X1 U13655 ( .B1(n842), .B2(n16864), .C1(n12715), .C2(n16858), .A(
        n13811), .ZN(n13808) );
  AOI22_X1 U13656 ( .A1(n16852), .A2(n8190), .B1(n16846), .B2(n8254), .ZN(
        n13811) );
  OAI221_X1 U13657 ( .B1(n841), .B2(n16864), .C1(n12714), .C2(n16858), .A(
        n13793), .ZN(n13790) );
  AOI22_X1 U13658 ( .A1(n16852), .A2(n8189), .B1(n16846), .B2(n8253), .ZN(
        n13793) );
  OAI221_X1 U13659 ( .B1(n7616), .B2(n16612), .C1(n7743), .C2(n16606), .A(
        n14985), .ZN(n14978) );
  AOI222_X1 U13660 ( .A1(n16600), .A2(n13382), .B1(n16594), .B2(n13190), .C1(
        n16588), .C2(n13062), .ZN(n14985) );
  OAI221_X1 U13661 ( .B1(n12998), .B2(n16511), .C1(n904), .C2(n16505), .A(
        n14993), .ZN(n14986) );
  AOI222_X1 U13662 ( .A1(n16499), .A2(n8892), .B1(n16493), .B2(n8764), .C1(
        n16487), .C2(n8828), .ZN(n14993) );
  OAI221_X1 U13663 ( .B1(n7614), .B2(n16612), .C1(n7741), .C2(n16606), .A(
        n14967), .ZN(n14960) );
  AOI222_X1 U13664 ( .A1(n16600), .A2(n13381), .B1(n16594), .B2(n13189), .C1(
        n16588), .C2(n13061), .ZN(n14967) );
  OAI221_X1 U13665 ( .B1(n12997), .B2(n16511), .C1(n903), .C2(n16505), .A(
        n14975), .ZN(n14968) );
  AOI222_X1 U13666 ( .A1(n16499), .A2(n8891), .B1(n16493), .B2(n8763), .C1(
        n16487), .C2(n8827), .ZN(n14975) );
  OAI221_X1 U13667 ( .B1(n7612), .B2(n16612), .C1(n7739), .C2(n16606), .A(
        n14949), .ZN(n14942) );
  AOI222_X1 U13668 ( .A1(n16600), .A2(n13380), .B1(n16594), .B2(n13188), .C1(
        n16588), .C2(n13060), .ZN(n14949) );
  OAI221_X1 U13669 ( .B1(n12996), .B2(n16511), .C1(n902), .C2(n16505), .A(
        n14957), .ZN(n14950) );
  AOI222_X1 U13670 ( .A1(n16499), .A2(n8890), .B1(n16493), .B2(n8762), .C1(
        n16487), .C2(n8826), .ZN(n14957) );
  OAI221_X1 U13671 ( .B1(n7610), .B2(n16612), .C1(n7737), .C2(n16606), .A(
        n14911), .ZN(n14890) );
  AOI222_X1 U13672 ( .A1(n16600), .A2(n13379), .B1(n16594), .B2(n13187), .C1(
        n16588), .C2(n13059), .ZN(n14911) );
  OAI221_X1 U13673 ( .B1(n12995), .B2(n16511), .C1(n901), .C2(n16505), .A(
        n14936), .ZN(n14915) );
  AOI222_X1 U13674 ( .A1(n16499), .A2(n8889), .B1(n16493), .B2(n8761), .C1(
        n16487), .C2(n8825), .ZN(n14936) );
  OAI221_X1 U13675 ( .B1(n7616), .B2(n16817), .C1(n7743), .C2(n16811), .A(
        n13777), .ZN(n13770) );
  AOI222_X1 U13676 ( .A1(n16805), .A2(n13382), .B1(n16799), .B2(n13190), .C1(
        n16793), .C2(n13062), .ZN(n13777) );
  OAI221_X1 U13677 ( .B1(n12998), .B2(n16716), .C1(n904), .C2(n16710), .A(
        n13785), .ZN(n13778) );
  AOI222_X1 U13678 ( .A1(n16704), .A2(n8892), .B1(n16698), .B2(n8764), .C1(
        n16692), .C2(n8828), .ZN(n13785) );
  OAI221_X1 U13679 ( .B1(n7614), .B2(n16817), .C1(n7741), .C2(n16811), .A(
        n13759), .ZN(n13752) );
  AOI222_X1 U13680 ( .A1(n16805), .A2(n13381), .B1(n16799), .B2(n13189), .C1(
        n16793), .C2(n13061), .ZN(n13759) );
  OAI221_X1 U13681 ( .B1(n12997), .B2(n16716), .C1(n903), .C2(n16710), .A(
        n13767), .ZN(n13760) );
  AOI222_X1 U13682 ( .A1(n16704), .A2(n8891), .B1(n16698), .B2(n8763), .C1(
        n16692), .C2(n8827), .ZN(n13767) );
  OAI221_X1 U13683 ( .B1(n7612), .B2(n16817), .C1(n7739), .C2(n16811), .A(
        n13741), .ZN(n13734) );
  AOI222_X1 U13684 ( .A1(n16805), .A2(n13380), .B1(n16799), .B2(n13188), .C1(
        n16793), .C2(n13060), .ZN(n13741) );
  OAI221_X1 U13685 ( .B1(n12996), .B2(n16716), .C1(n902), .C2(n16710), .A(
        n13749), .ZN(n13742) );
  AOI222_X1 U13686 ( .A1(n16704), .A2(n8890), .B1(n16698), .B2(n8762), .C1(
        n16692), .C2(n8826), .ZN(n13749) );
  OAI221_X1 U13687 ( .B1(n7610), .B2(n16817), .C1(n7737), .C2(n16811), .A(
        n13703), .ZN(n13682) );
  AOI222_X1 U13688 ( .A1(n16805), .A2(n13379), .B1(n16799), .B2(n13187), .C1(
        n16793), .C2(n13059), .ZN(n13703) );
  OAI221_X1 U13689 ( .B1(n12995), .B2(n16716), .C1(n901), .C2(n16710), .A(
        n13728), .ZN(n13707) );
  AOI222_X1 U13690 ( .A1(n16704), .A2(n8889), .B1(n16698), .B2(n8761), .C1(
        n16692), .C2(n8825), .ZN(n13728) );
  OAI221_X1 U13691 ( .B1(n13477), .B2(n16737), .C1(n999), .C2(n16731), .A(
        n14342), .ZN(n14337) );
  AOI22_X1 U13692 ( .A1(n16725), .A2(n12232), .B1(n16719), .B2(n12424), .ZN(
        n14342) );
  OAI221_X1 U13693 ( .B1(n13476), .B2(n16737), .C1(n998), .C2(n16731), .A(
        n14324), .ZN(n14319) );
  AOI22_X1 U13694 ( .A1(n16725), .A2(n12231), .B1(n16719), .B2(n12423), .ZN(
        n14324) );
  OAI221_X1 U13695 ( .B1(n13475), .B2(n16737), .C1(n997), .C2(n16731), .A(
        n14306), .ZN(n14301) );
  AOI22_X1 U13696 ( .A1(n16725), .A2(n12230), .B1(n16719), .B2(n12422), .ZN(
        n14306) );
  OAI221_X1 U13697 ( .B1(n13474), .B2(n16737), .C1(n996), .C2(n16731), .A(
        n14288), .ZN(n14283) );
  AOI22_X1 U13698 ( .A1(n16725), .A2(n12229), .B1(n16719), .B2(n12421), .ZN(
        n14288) );
  OAI221_X1 U13699 ( .B1(n13473), .B2(n16737), .C1(n995), .C2(n16731), .A(
        n14270), .ZN(n14265) );
  AOI22_X1 U13700 ( .A1(n16725), .A2(n12228), .B1(n16719), .B2(n12420), .ZN(
        n14270) );
  OAI221_X1 U13701 ( .B1(n13472), .B2(n16737), .C1(n994), .C2(n16731), .A(
        n14252), .ZN(n14247) );
  AOI22_X1 U13702 ( .A1(n16725), .A2(n12227), .B1(n16719), .B2(n12419), .ZN(
        n14252) );
  OAI221_X1 U13703 ( .B1(n13471), .B2(n16737), .C1(n993), .C2(n16731), .A(
        n14234), .ZN(n14229) );
  AOI22_X1 U13704 ( .A1(n16725), .A2(n12226), .B1(n16719), .B2(n12418), .ZN(
        n14234) );
  OAI221_X1 U13705 ( .B1(n13470), .B2(n16738), .C1(n992), .C2(n16732), .A(
        n14216), .ZN(n14211) );
  AOI22_X1 U13706 ( .A1(n16726), .A2(n12225), .B1(n16720), .B2(n12417), .ZN(
        n14216) );
  OAI221_X1 U13707 ( .B1(n13469), .B2(n16738), .C1(n991), .C2(n16732), .A(
        n14198), .ZN(n14193) );
  AOI22_X1 U13708 ( .A1(n16726), .A2(n12224), .B1(n16720), .B2(n12416), .ZN(
        n14198) );
  OAI221_X1 U13709 ( .B1(n13468), .B2(n16738), .C1(n990), .C2(n16732), .A(
        n14180), .ZN(n14175) );
  AOI22_X1 U13710 ( .A1(n16726), .A2(n12223), .B1(n16720), .B2(n12415), .ZN(
        n14180) );
  OAI221_X1 U13711 ( .B1(n13467), .B2(n16738), .C1(n989), .C2(n16732), .A(
        n14162), .ZN(n14157) );
  AOI22_X1 U13712 ( .A1(n16726), .A2(n12222), .B1(n16720), .B2(n12414), .ZN(
        n14162) );
  OAI221_X1 U13713 ( .B1(n13466), .B2(n16738), .C1(n988), .C2(n16732), .A(
        n14144), .ZN(n14139) );
  AOI22_X1 U13714 ( .A1(n16726), .A2(n12221), .B1(n16720), .B2(n12413), .ZN(
        n14144) );
  OAI221_X1 U13715 ( .B1(n13465), .B2(n16738), .C1(n987), .C2(n16732), .A(
        n14126), .ZN(n14121) );
  AOI22_X1 U13716 ( .A1(n16726), .A2(n12220), .B1(n16720), .B2(n12412), .ZN(
        n14126) );
  OAI221_X1 U13717 ( .B1(n13464), .B2(n16738), .C1(n986), .C2(n16732), .A(
        n14108), .ZN(n14103) );
  AOI22_X1 U13718 ( .A1(n16726), .A2(n12219), .B1(n16720), .B2(n12411), .ZN(
        n14108) );
  OAI221_X1 U13719 ( .B1(n13463), .B2(n16738), .C1(n985), .C2(n16732), .A(
        n14090), .ZN(n14085) );
  AOI22_X1 U13720 ( .A1(n16726), .A2(n12218), .B1(n16720), .B2(n12410), .ZN(
        n14090) );
  OAI221_X1 U13721 ( .B1(n13462), .B2(n16738), .C1(n984), .C2(n16732), .A(
        n14072), .ZN(n14067) );
  AOI22_X1 U13722 ( .A1(n16726), .A2(n12217), .B1(n16720), .B2(n12409), .ZN(
        n14072) );
  OAI221_X1 U13723 ( .B1(n13461), .B2(n16738), .C1(n983), .C2(n16732), .A(
        n14054), .ZN(n14049) );
  AOI22_X1 U13724 ( .A1(n16726), .A2(n12216), .B1(n16720), .B2(n12408), .ZN(
        n14054) );
  OAI221_X1 U13725 ( .B1(n13460), .B2(n16738), .C1(n982), .C2(n16732), .A(
        n14036), .ZN(n14031) );
  AOI22_X1 U13726 ( .A1(n16726), .A2(n12215), .B1(n16720), .B2(n12407), .ZN(
        n14036) );
  OAI221_X1 U13727 ( .B1(n13459), .B2(n16738), .C1(n981), .C2(n16732), .A(
        n14018), .ZN(n14013) );
  AOI22_X1 U13728 ( .A1(n16726), .A2(n12214), .B1(n16720), .B2(n12406), .ZN(
        n14018) );
  OAI221_X1 U13729 ( .B1(n7736), .B2(n16607), .C1(n7863), .C2(n16601), .A(
        n16076), .ZN(n16058) );
  AOI222_X1 U13730 ( .A1(n16595), .A2(n13442), .B1(n16589), .B2(n13250), .C1(
        n16583), .C2(n13122), .ZN(n16076) );
  OAI221_X1 U13731 ( .B1(n7734), .B2(n16607), .C1(n7861), .C2(n16601), .A(
        n16047), .ZN(n16040) );
  AOI222_X1 U13732 ( .A1(n16595), .A2(n13441), .B1(n16589), .B2(n13249), .C1(
        n16583), .C2(n13121), .ZN(n16047) );
  OAI221_X1 U13733 ( .B1(n7732), .B2(n16607), .C1(n7859), .C2(n16601), .A(
        n16029), .ZN(n16022) );
  AOI222_X1 U13734 ( .A1(n16595), .A2(n13440), .B1(n16589), .B2(n13248), .C1(
        n16583), .C2(n13120), .ZN(n16029) );
  OAI221_X1 U13735 ( .B1(n7730), .B2(n16607), .C1(n7857), .C2(n16601), .A(
        n16011), .ZN(n16004) );
  AOI222_X1 U13736 ( .A1(n16595), .A2(n13439), .B1(n16589), .B2(n13247), .C1(
        n16583), .C2(n13119), .ZN(n16011) );
  OAI221_X1 U13737 ( .B1(n7728), .B2(n16607), .C1(n7855), .C2(n16601), .A(
        n15993), .ZN(n15986) );
  AOI222_X1 U13738 ( .A1(n16595), .A2(n13438), .B1(n16589), .B2(n13246), .C1(
        n16583), .C2(n13118), .ZN(n15993) );
  OAI221_X1 U13739 ( .B1(n7726), .B2(n16607), .C1(n7853), .C2(n16601), .A(
        n15975), .ZN(n15968) );
  AOI222_X1 U13740 ( .A1(n16595), .A2(n13437), .B1(n16589), .B2(n13245), .C1(
        n16583), .C2(n13117), .ZN(n15975) );
  OAI221_X1 U13741 ( .B1(n7724), .B2(n16607), .C1(n7851), .C2(n16601), .A(
        n15957), .ZN(n15950) );
  AOI222_X1 U13742 ( .A1(n16595), .A2(n13436), .B1(n16589), .B2(n13244), .C1(
        n16583), .C2(n13116), .ZN(n15957) );
  OAI221_X1 U13743 ( .B1(n7722), .B2(n16607), .C1(n7849), .C2(n16601), .A(
        n15939), .ZN(n15932) );
  AOI222_X1 U13744 ( .A1(n16595), .A2(n13435), .B1(n16589), .B2(n13243), .C1(
        n16583), .C2(n13115), .ZN(n15939) );
  OAI221_X1 U13745 ( .B1(n7720), .B2(n16607), .C1(n7847), .C2(n16601), .A(
        n15921), .ZN(n15914) );
  AOI222_X1 U13746 ( .A1(n16595), .A2(n13434), .B1(n16589), .B2(n13242), .C1(
        n16583), .C2(n13114), .ZN(n15921) );
  OAI221_X1 U13747 ( .B1(n7718), .B2(n16607), .C1(n7845), .C2(n16601), .A(
        n15903), .ZN(n15896) );
  AOI222_X1 U13748 ( .A1(n16595), .A2(n13433), .B1(n16589), .B2(n13241), .C1(
        n16583), .C2(n13113), .ZN(n15903) );
  OAI221_X1 U13749 ( .B1(n7716), .B2(n16607), .C1(n7843), .C2(n16601), .A(
        n15885), .ZN(n15878) );
  AOI222_X1 U13750 ( .A1(n16595), .A2(n13432), .B1(n16589), .B2(n13240), .C1(
        n16583), .C2(n13112), .ZN(n15885) );
  OAI221_X1 U13751 ( .B1(n7714), .B2(n16607), .C1(n7841), .C2(n16601), .A(
        n15867), .ZN(n15860) );
  AOI222_X1 U13752 ( .A1(n16595), .A2(n13431), .B1(n16589), .B2(n13239), .C1(
        n16583), .C2(n13111), .ZN(n15867) );
  OAI221_X1 U13753 ( .B1(n7712), .B2(n16608), .C1(n7839), .C2(n16602), .A(
        n15849), .ZN(n15842) );
  AOI222_X1 U13754 ( .A1(n16596), .A2(n13430), .B1(n16590), .B2(n13238), .C1(
        n16584), .C2(n13110), .ZN(n15849) );
  OAI221_X1 U13755 ( .B1(n7710), .B2(n16608), .C1(n7837), .C2(n16602), .A(
        n15831), .ZN(n15824) );
  AOI222_X1 U13756 ( .A1(n16596), .A2(n13429), .B1(n16590), .B2(n13237), .C1(
        n16584), .C2(n13109), .ZN(n15831) );
  OAI221_X1 U13757 ( .B1(n7708), .B2(n16608), .C1(n7835), .C2(n16602), .A(
        n15813), .ZN(n15806) );
  AOI222_X1 U13758 ( .A1(n16596), .A2(n13428), .B1(n16590), .B2(n13236), .C1(
        n16584), .C2(n13108), .ZN(n15813) );
  OAI221_X1 U13759 ( .B1(n7706), .B2(n16608), .C1(n7833), .C2(n16602), .A(
        n15795), .ZN(n15788) );
  AOI222_X1 U13760 ( .A1(n16596), .A2(n13427), .B1(n16590), .B2(n13235), .C1(
        n16584), .C2(n13107), .ZN(n15795) );
  OAI221_X1 U13761 ( .B1(n7704), .B2(n16608), .C1(n7831), .C2(n16602), .A(
        n15777), .ZN(n15770) );
  AOI222_X1 U13762 ( .A1(n16596), .A2(n13426), .B1(n16590), .B2(n13234), .C1(
        n16584), .C2(n13106), .ZN(n15777) );
  OAI221_X1 U13763 ( .B1(n7702), .B2(n16608), .C1(n7829), .C2(n16602), .A(
        n15759), .ZN(n15752) );
  AOI222_X1 U13764 ( .A1(n16596), .A2(n13425), .B1(n16590), .B2(n13233), .C1(
        n16584), .C2(n13105), .ZN(n15759) );
  OAI221_X1 U13765 ( .B1(n7700), .B2(n16608), .C1(n7827), .C2(n16602), .A(
        n15741), .ZN(n15734) );
  AOI222_X1 U13766 ( .A1(n16596), .A2(n13424), .B1(n16590), .B2(n13232), .C1(
        n16584), .C2(n13104), .ZN(n15741) );
  OAI221_X1 U13767 ( .B1(n7698), .B2(n16608), .C1(n7825), .C2(n16602), .A(
        n15723), .ZN(n15716) );
  AOI222_X1 U13768 ( .A1(n16596), .A2(n13423), .B1(n16590), .B2(n13231), .C1(
        n16584), .C2(n13103), .ZN(n15723) );
  OAI221_X1 U13769 ( .B1(n7696), .B2(n16608), .C1(n7823), .C2(n16602), .A(
        n15705), .ZN(n15698) );
  AOI222_X1 U13770 ( .A1(n16596), .A2(n13422), .B1(n16590), .B2(n13230), .C1(
        n16584), .C2(n13102), .ZN(n15705) );
  OAI221_X1 U13771 ( .B1(n7694), .B2(n16608), .C1(n7821), .C2(n16602), .A(
        n15687), .ZN(n15680) );
  AOI222_X1 U13772 ( .A1(n16596), .A2(n13421), .B1(n16590), .B2(n13229), .C1(
        n16584), .C2(n13101), .ZN(n15687) );
  OAI221_X1 U13773 ( .B1(n7692), .B2(n16608), .C1(n7819), .C2(n16602), .A(
        n15669), .ZN(n15662) );
  AOI222_X1 U13774 ( .A1(n16596), .A2(n13420), .B1(n16590), .B2(n13228), .C1(
        n16584), .C2(n13100), .ZN(n15669) );
  OAI221_X1 U13775 ( .B1(n7690), .B2(n16608), .C1(n7817), .C2(n16602), .A(
        n15651), .ZN(n15644) );
  AOI222_X1 U13776 ( .A1(n16596), .A2(n13419), .B1(n16590), .B2(n13227), .C1(
        n16584), .C2(n13099), .ZN(n15651) );
  OAI221_X1 U13777 ( .B1(n7688), .B2(n16609), .C1(n7815), .C2(n16603), .A(
        n15633), .ZN(n15626) );
  AOI222_X1 U13778 ( .A1(n16597), .A2(n13418), .B1(n16591), .B2(n13226), .C1(
        n16585), .C2(n13098), .ZN(n15633) );
  OAI221_X1 U13779 ( .B1(n7686), .B2(n16609), .C1(n7813), .C2(n16603), .A(
        n15615), .ZN(n15608) );
  AOI222_X1 U13780 ( .A1(n16597), .A2(n13417), .B1(n16591), .B2(n13225), .C1(
        n16585), .C2(n13097), .ZN(n15615) );
  OAI221_X1 U13781 ( .B1(n7684), .B2(n16609), .C1(n7811), .C2(n16603), .A(
        n15597), .ZN(n15590) );
  AOI222_X1 U13782 ( .A1(n16597), .A2(n13416), .B1(n16591), .B2(n13224), .C1(
        n16585), .C2(n13096), .ZN(n15597) );
  OAI221_X1 U13783 ( .B1(n7682), .B2(n16609), .C1(n7809), .C2(n16603), .A(
        n15579), .ZN(n15572) );
  AOI222_X1 U13784 ( .A1(n16597), .A2(n13415), .B1(n16591), .B2(n13223), .C1(
        n16585), .C2(n13095), .ZN(n15579) );
  OAI221_X1 U13785 ( .B1(n7680), .B2(n16609), .C1(n7807), .C2(n16603), .A(
        n15561), .ZN(n15554) );
  AOI222_X1 U13786 ( .A1(n16597), .A2(n13414), .B1(n16591), .B2(n13222), .C1(
        n16585), .C2(n13094), .ZN(n15561) );
  OAI221_X1 U13787 ( .B1(n7678), .B2(n16609), .C1(n7805), .C2(n16603), .A(
        n15543), .ZN(n15536) );
  AOI222_X1 U13788 ( .A1(n16597), .A2(n13413), .B1(n16591), .B2(n13221), .C1(
        n16585), .C2(n13093), .ZN(n15543) );
  OAI221_X1 U13789 ( .B1(n7676), .B2(n16609), .C1(n7803), .C2(n16603), .A(
        n15525), .ZN(n15518) );
  AOI222_X1 U13790 ( .A1(n16597), .A2(n13412), .B1(n16591), .B2(n13220), .C1(
        n16585), .C2(n13092), .ZN(n15525) );
  OAI221_X1 U13791 ( .B1(n7674), .B2(n16609), .C1(n7801), .C2(n16603), .A(
        n15507), .ZN(n15500) );
  AOI222_X1 U13792 ( .A1(n16597), .A2(n13411), .B1(n16591), .B2(n13219), .C1(
        n16585), .C2(n13091), .ZN(n15507) );
  OAI221_X1 U13793 ( .B1(n7672), .B2(n16609), .C1(n7799), .C2(n16603), .A(
        n15489), .ZN(n15482) );
  AOI222_X1 U13794 ( .A1(n16597), .A2(n13410), .B1(n16591), .B2(n13218), .C1(
        n16585), .C2(n13090), .ZN(n15489) );
  OAI221_X1 U13795 ( .B1(n7670), .B2(n16609), .C1(n7797), .C2(n16603), .A(
        n15471), .ZN(n15464) );
  AOI222_X1 U13796 ( .A1(n16597), .A2(n13409), .B1(n16591), .B2(n13217), .C1(
        n16585), .C2(n13089), .ZN(n15471) );
  OAI221_X1 U13797 ( .B1(n7668), .B2(n16609), .C1(n7795), .C2(n16603), .A(
        n15453), .ZN(n15446) );
  AOI222_X1 U13798 ( .A1(n16597), .A2(n13408), .B1(n16591), .B2(n13216), .C1(
        n16585), .C2(n13088), .ZN(n15453) );
  OAI221_X1 U13799 ( .B1(n7666), .B2(n16609), .C1(n7793), .C2(n16603), .A(
        n15435), .ZN(n15428) );
  AOI222_X1 U13800 ( .A1(n16597), .A2(n13407), .B1(n16591), .B2(n13215), .C1(
        n16585), .C2(n13087), .ZN(n15435) );
  OAI221_X1 U13801 ( .B1(n7664), .B2(n16610), .C1(n7791), .C2(n16604), .A(
        n15417), .ZN(n15410) );
  AOI222_X1 U13802 ( .A1(n16598), .A2(n13406), .B1(n16592), .B2(n13214), .C1(
        n16586), .C2(n13086), .ZN(n15417) );
  OAI221_X1 U13803 ( .B1(n7662), .B2(n16610), .C1(n7789), .C2(n16604), .A(
        n15399), .ZN(n15392) );
  AOI222_X1 U13804 ( .A1(n16598), .A2(n13405), .B1(n16592), .B2(n13213), .C1(
        n16586), .C2(n13085), .ZN(n15399) );
  OAI221_X1 U13805 ( .B1(n7660), .B2(n16610), .C1(n7787), .C2(n16604), .A(
        n15381), .ZN(n15374) );
  AOI222_X1 U13806 ( .A1(n16598), .A2(n13404), .B1(n16592), .B2(n13212), .C1(
        n16586), .C2(n13084), .ZN(n15381) );
  OAI221_X1 U13807 ( .B1(n7658), .B2(n16610), .C1(n7785), .C2(n16604), .A(
        n15363), .ZN(n15356) );
  AOI222_X1 U13808 ( .A1(n16598), .A2(n13403), .B1(n16592), .B2(n13211), .C1(
        n16586), .C2(n13083), .ZN(n15363) );
  OAI221_X1 U13809 ( .B1(n7656), .B2(n16610), .C1(n7783), .C2(n16604), .A(
        n15345), .ZN(n15338) );
  AOI222_X1 U13810 ( .A1(n16598), .A2(n13402), .B1(n16592), .B2(n13210), .C1(
        n16586), .C2(n13082), .ZN(n15345) );
  OAI221_X1 U13811 ( .B1(n7654), .B2(n16610), .C1(n7781), .C2(n16604), .A(
        n15327), .ZN(n15320) );
  AOI222_X1 U13812 ( .A1(n16598), .A2(n13401), .B1(n16592), .B2(n13209), .C1(
        n16586), .C2(n13081), .ZN(n15327) );
  OAI221_X1 U13813 ( .B1(n7652), .B2(n16610), .C1(n7779), .C2(n16604), .A(
        n15309), .ZN(n15302) );
  AOI222_X1 U13814 ( .A1(n16598), .A2(n13400), .B1(n16592), .B2(n13208), .C1(
        n16586), .C2(n13080), .ZN(n15309) );
  OAI221_X1 U13815 ( .B1(n7650), .B2(n16610), .C1(n7777), .C2(n16604), .A(
        n15291), .ZN(n15284) );
  AOI222_X1 U13816 ( .A1(n16598), .A2(n13399), .B1(n16592), .B2(n13207), .C1(
        n16586), .C2(n13079), .ZN(n15291) );
  OAI221_X1 U13817 ( .B1(n7648), .B2(n16610), .C1(n7775), .C2(n16604), .A(
        n15273), .ZN(n15266) );
  AOI222_X1 U13818 ( .A1(n16598), .A2(n13398), .B1(n16592), .B2(n13206), .C1(
        n16586), .C2(n13078), .ZN(n15273) );
  OAI221_X1 U13819 ( .B1(n7646), .B2(n16610), .C1(n7773), .C2(n16604), .A(
        n15255), .ZN(n15248) );
  AOI222_X1 U13820 ( .A1(n16598), .A2(n13397), .B1(n16592), .B2(n13205), .C1(
        n16586), .C2(n13077), .ZN(n15255) );
  OAI221_X1 U13821 ( .B1(n7644), .B2(n16610), .C1(n7771), .C2(n16604), .A(
        n15237), .ZN(n15230) );
  AOI222_X1 U13822 ( .A1(n16598), .A2(n13396), .B1(n16592), .B2(n13204), .C1(
        n16586), .C2(n13076), .ZN(n15237) );
  OAI221_X1 U13823 ( .B1(n7642), .B2(n16610), .C1(n7769), .C2(n16604), .A(
        n15219), .ZN(n15212) );
  AOI222_X1 U13824 ( .A1(n16598), .A2(n13395), .B1(n16592), .B2(n13203), .C1(
        n16586), .C2(n13075), .ZN(n15219) );
  OAI221_X1 U13825 ( .B1(n7640), .B2(n16611), .C1(n7767), .C2(n16605), .A(
        n15201), .ZN(n15194) );
  AOI222_X1 U13826 ( .A1(n16599), .A2(n13394), .B1(n16593), .B2(n13202), .C1(
        n16587), .C2(n13074), .ZN(n15201) );
  OAI221_X1 U13827 ( .B1(n7638), .B2(n16611), .C1(n7765), .C2(n16605), .A(
        n15183), .ZN(n15176) );
  AOI222_X1 U13828 ( .A1(n16599), .A2(n13393), .B1(n16593), .B2(n13201), .C1(
        n16587), .C2(n13073), .ZN(n15183) );
  OAI221_X1 U13829 ( .B1(n7636), .B2(n16611), .C1(n7763), .C2(n16605), .A(
        n15165), .ZN(n15158) );
  AOI222_X1 U13830 ( .A1(n16599), .A2(n13392), .B1(n16593), .B2(n13200), .C1(
        n16587), .C2(n13072), .ZN(n15165) );
  OAI221_X1 U13831 ( .B1(n7634), .B2(n16611), .C1(n7761), .C2(n16605), .A(
        n15147), .ZN(n15140) );
  AOI222_X1 U13832 ( .A1(n16599), .A2(n13391), .B1(n16593), .B2(n13199), .C1(
        n16587), .C2(n13071), .ZN(n15147) );
  OAI221_X1 U13833 ( .B1(n7632), .B2(n16611), .C1(n7759), .C2(n16605), .A(
        n15129), .ZN(n15122) );
  AOI222_X1 U13834 ( .A1(n16599), .A2(n13390), .B1(n16593), .B2(n13198), .C1(
        n16587), .C2(n13070), .ZN(n15129) );
  OAI221_X1 U13835 ( .B1(n7630), .B2(n16611), .C1(n7757), .C2(n16605), .A(
        n15111), .ZN(n15104) );
  AOI222_X1 U13836 ( .A1(n16599), .A2(n13389), .B1(n16593), .B2(n13197), .C1(
        n16587), .C2(n13069), .ZN(n15111) );
  OAI221_X1 U13837 ( .B1(n7628), .B2(n16611), .C1(n7755), .C2(n16605), .A(
        n15093), .ZN(n15086) );
  AOI222_X1 U13838 ( .A1(n16599), .A2(n13388), .B1(n16593), .B2(n13196), .C1(
        n16587), .C2(n13068), .ZN(n15093) );
  OAI221_X1 U13839 ( .B1(n7626), .B2(n16611), .C1(n7753), .C2(n16605), .A(
        n15075), .ZN(n15068) );
  AOI222_X1 U13840 ( .A1(n16599), .A2(n13387), .B1(n16593), .B2(n13195), .C1(
        n16587), .C2(n13067), .ZN(n15075) );
  OAI221_X1 U13841 ( .B1(n7624), .B2(n16611), .C1(n7751), .C2(n16605), .A(
        n15057), .ZN(n15050) );
  AOI222_X1 U13842 ( .A1(n16599), .A2(n13386), .B1(n16593), .B2(n13194), .C1(
        n16587), .C2(n13066), .ZN(n15057) );
  OAI221_X1 U13843 ( .B1(n7622), .B2(n16611), .C1(n7749), .C2(n16605), .A(
        n15039), .ZN(n15032) );
  AOI222_X1 U13844 ( .A1(n16599), .A2(n13385), .B1(n16593), .B2(n13193), .C1(
        n16587), .C2(n13065), .ZN(n15039) );
  OAI221_X1 U13845 ( .B1(n7620), .B2(n16611), .C1(n7747), .C2(n16605), .A(
        n15021), .ZN(n15014) );
  AOI222_X1 U13846 ( .A1(n16599), .A2(n13384), .B1(n16593), .B2(n13192), .C1(
        n16587), .C2(n13064), .ZN(n15021) );
  OAI221_X1 U13847 ( .B1(n7618), .B2(n16611), .C1(n7745), .C2(n16605), .A(
        n15003), .ZN(n14996) );
  AOI222_X1 U13848 ( .A1(n16599), .A2(n13383), .B1(n16593), .B2(n13191), .C1(
        n16587), .C2(n13063), .ZN(n15003) );
  OAI221_X1 U13849 ( .B1(n7736), .B2(n16812), .C1(n7863), .C2(n16806), .A(
        n14868), .ZN(n14850) );
  AOI222_X1 U13850 ( .A1(n16800), .A2(n13442), .B1(n16794), .B2(n13250), .C1(
        n16788), .C2(n13122), .ZN(n14868) );
  OAI221_X1 U13851 ( .B1(n7734), .B2(n16812), .C1(n7861), .C2(n16806), .A(
        n14839), .ZN(n14832) );
  AOI222_X1 U13852 ( .A1(n16800), .A2(n13441), .B1(n16794), .B2(n13249), .C1(
        n16788), .C2(n13121), .ZN(n14839) );
  OAI221_X1 U13853 ( .B1(n7732), .B2(n16812), .C1(n7859), .C2(n16806), .A(
        n14821), .ZN(n14814) );
  AOI222_X1 U13854 ( .A1(n16800), .A2(n13440), .B1(n16794), .B2(n13248), .C1(
        n16788), .C2(n13120), .ZN(n14821) );
  OAI221_X1 U13855 ( .B1(n7730), .B2(n16812), .C1(n7857), .C2(n16806), .A(
        n14803), .ZN(n14796) );
  AOI222_X1 U13856 ( .A1(n16800), .A2(n13439), .B1(n16794), .B2(n13247), .C1(
        n16788), .C2(n13119), .ZN(n14803) );
  OAI221_X1 U13857 ( .B1(n7728), .B2(n16812), .C1(n7855), .C2(n16806), .A(
        n14785), .ZN(n14778) );
  AOI222_X1 U13858 ( .A1(n16800), .A2(n13438), .B1(n16794), .B2(n13246), .C1(
        n16788), .C2(n13118), .ZN(n14785) );
  OAI221_X1 U13859 ( .B1(n7726), .B2(n16812), .C1(n7853), .C2(n16806), .A(
        n14767), .ZN(n14760) );
  AOI222_X1 U13860 ( .A1(n16800), .A2(n13437), .B1(n16794), .B2(n13245), .C1(
        n16788), .C2(n13117), .ZN(n14767) );
  OAI221_X1 U13861 ( .B1(n7724), .B2(n16812), .C1(n7851), .C2(n16806), .A(
        n14749), .ZN(n14742) );
  AOI222_X1 U13862 ( .A1(n16800), .A2(n13436), .B1(n16794), .B2(n13244), .C1(
        n16788), .C2(n13116), .ZN(n14749) );
  OAI221_X1 U13863 ( .B1(n7722), .B2(n16812), .C1(n7849), .C2(n16806), .A(
        n14731), .ZN(n14724) );
  AOI222_X1 U13864 ( .A1(n16800), .A2(n13435), .B1(n16794), .B2(n13243), .C1(
        n16788), .C2(n13115), .ZN(n14731) );
  OAI221_X1 U13865 ( .B1(n7720), .B2(n16812), .C1(n7847), .C2(n16806), .A(
        n14713), .ZN(n14706) );
  AOI222_X1 U13866 ( .A1(n16800), .A2(n13434), .B1(n16794), .B2(n13242), .C1(
        n16788), .C2(n13114), .ZN(n14713) );
  OAI221_X1 U13867 ( .B1(n7718), .B2(n16812), .C1(n7845), .C2(n16806), .A(
        n14695), .ZN(n14688) );
  AOI222_X1 U13868 ( .A1(n16800), .A2(n13433), .B1(n16794), .B2(n13241), .C1(
        n16788), .C2(n13113), .ZN(n14695) );
  OAI221_X1 U13869 ( .B1(n7716), .B2(n16812), .C1(n7843), .C2(n16806), .A(
        n14677), .ZN(n14670) );
  AOI222_X1 U13870 ( .A1(n16800), .A2(n13432), .B1(n16794), .B2(n13240), .C1(
        n16788), .C2(n13112), .ZN(n14677) );
  OAI221_X1 U13871 ( .B1(n7714), .B2(n16812), .C1(n7841), .C2(n16806), .A(
        n14659), .ZN(n14652) );
  AOI222_X1 U13872 ( .A1(n16800), .A2(n13431), .B1(n16794), .B2(n13239), .C1(
        n16788), .C2(n13111), .ZN(n14659) );
  OAI221_X1 U13873 ( .B1(n7712), .B2(n16813), .C1(n7839), .C2(n16807), .A(
        n14641), .ZN(n14634) );
  AOI222_X1 U13874 ( .A1(n16801), .A2(n13430), .B1(n16795), .B2(n13238), .C1(
        n16789), .C2(n13110), .ZN(n14641) );
  OAI221_X1 U13875 ( .B1(n7710), .B2(n16813), .C1(n7837), .C2(n16807), .A(
        n14623), .ZN(n14616) );
  AOI222_X1 U13876 ( .A1(n16801), .A2(n13429), .B1(n16795), .B2(n13237), .C1(
        n16789), .C2(n13109), .ZN(n14623) );
  OAI221_X1 U13877 ( .B1(n7708), .B2(n16813), .C1(n7835), .C2(n16807), .A(
        n14605), .ZN(n14598) );
  AOI222_X1 U13878 ( .A1(n16801), .A2(n13428), .B1(n16795), .B2(n13236), .C1(
        n16789), .C2(n13108), .ZN(n14605) );
  OAI221_X1 U13879 ( .B1(n7706), .B2(n16813), .C1(n7833), .C2(n16807), .A(
        n14587), .ZN(n14580) );
  AOI222_X1 U13880 ( .A1(n16801), .A2(n13427), .B1(n16795), .B2(n13235), .C1(
        n16789), .C2(n13107), .ZN(n14587) );
  OAI221_X1 U13881 ( .B1(n7704), .B2(n16813), .C1(n7831), .C2(n16807), .A(
        n14569), .ZN(n14562) );
  AOI222_X1 U13882 ( .A1(n16801), .A2(n13426), .B1(n16795), .B2(n13234), .C1(
        n16789), .C2(n13106), .ZN(n14569) );
  OAI221_X1 U13883 ( .B1(n7702), .B2(n16813), .C1(n7829), .C2(n16807), .A(
        n14551), .ZN(n14544) );
  AOI222_X1 U13884 ( .A1(n16801), .A2(n13425), .B1(n16795), .B2(n13233), .C1(
        n16789), .C2(n13105), .ZN(n14551) );
  OAI221_X1 U13885 ( .B1(n7700), .B2(n16813), .C1(n7827), .C2(n16807), .A(
        n14533), .ZN(n14526) );
  AOI222_X1 U13886 ( .A1(n16801), .A2(n13424), .B1(n16795), .B2(n13232), .C1(
        n16789), .C2(n13104), .ZN(n14533) );
  OAI221_X1 U13887 ( .B1(n7698), .B2(n16813), .C1(n7825), .C2(n16807), .A(
        n14515), .ZN(n14508) );
  AOI222_X1 U13888 ( .A1(n16801), .A2(n13423), .B1(n16795), .B2(n13231), .C1(
        n16789), .C2(n13103), .ZN(n14515) );
  OAI221_X1 U13889 ( .B1(n7696), .B2(n16813), .C1(n7823), .C2(n16807), .A(
        n14497), .ZN(n14490) );
  AOI222_X1 U13890 ( .A1(n16801), .A2(n13422), .B1(n16795), .B2(n13230), .C1(
        n16789), .C2(n13102), .ZN(n14497) );
  OAI221_X1 U13891 ( .B1(n7694), .B2(n16813), .C1(n7821), .C2(n16807), .A(
        n14479), .ZN(n14472) );
  AOI222_X1 U13892 ( .A1(n16801), .A2(n13421), .B1(n16795), .B2(n13229), .C1(
        n16789), .C2(n13101), .ZN(n14479) );
  OAI221_X1 U13893 ( .B1(n7692), .B2(n16813), .C1(n7819), .C2(n16807), .A(
        n14461), .ZN(n14454) );
  AOI222_X1 U13894 ( .A1(n16801), .A2(n13420), .B1(n16795), .B2(n13228), .C1(
        n16789), .C2(n13100), .ZN(n14461) );
  OAI221_X1 U13895 ( .B1(n7690), .B2(n16813), .C1(n7817), .C2(n16807), .A(
        n14443), .ZN(n14436) );
  AOI222_X1 U13896 ( .A1(n16801), .A2(n13419), .B1(n16795), .B2(n13227), .C1(
        n16789), .C2(n13099), .ZN(n14443) );
  OAI221_X1 U13897 ( .B1(n7688), .B2(n16814), .C1(n7815), .C2(n16808), .A(
        n14425), .ZN(n14418) );
  AOI222_X1 U13898 ( .A1(n16802), .A2(n13418), .B1(n16796), .B2(n13226), .C1(
        n16790), .C2(n13098), .ZN(n14425) );
  OAI221_X1 U13899 ( .B1(n7686), .B2(n16814), .C1(n7813), .C2(n16808), .A(
        n14407), .ZN(n14400) );
  AOI222_X1 U13900 ( .A1(n16802), .A2(n13417), .B1(n16796), .B2(n13225), .C1(
        n16790), .C2(n13097), .ZN(n14407) );
  OAI221_X1 U13901 ( .B1(n7684), .B2(n16814), .C1(n7811), .C2(n16808), .A(
        n14389), .ZN(n14382) );
  AOI222_X1 U13902 ( .A1(n16802), .A2(n13416), .B1(n16796), .B2(n13224), .C1(
        n16790), .C2(n13096), .ZN(n14389) );
  OAI221_X1 U13903 ( .B1(n7682), .B2(n16814), .C1(n7809), .C2(n16808), .A(
        n14371), .ZN(n14364) );
  AOI222_X1 U13904 ( .A1(n16802), .A2(n13415), .B1(n16796), .B2(n13223), .C1(
        n16790), .C2(n13095), .ZN(n14371) );
  OAI221_X1 U13905 ( .B1(n7680), .B2(n16814), .C1(n7807), .C2(n16808), .A(
        n14353), .ZN(n14346) );
  AOI222_X1 U13906 ( .A1(n16802), .A2(n13414), .B1(n16796), .B2(n13222), .C1(
        n16790), .C2(n13094), .ZN(n14353) );
  OAI221_X1 U13907 ( .B1(n7678), .B2(n16814), .C1(n7805), .C2(n16808), .A(
        n14335), .ZN(n14328) );
  AOI222_X1 U13908 ( .A1(n16802), .A2(n13413), .B1(n16796), .B2(n13221), .C1(
        n16790), .C2(n13093), .ZN(n14335) );
  OAI221_X1 U13909 ( .B1(n7676), .B2(n16814), .C1(n7803), .C2(n16808), .A(
        n14317), .ZN(n14310) );
  AOI222_X1 U13910 ( .A1(n16802), .A2(n13412), .B1(n16796), .B2(n13220), .C1(
        n16790), .C2(n13092), .ZN(n14317) );
  OAI221_X1 U13911 ( .B1(n7674), .B2(n16814), .C1(n7801), .C2(n16808), .A(
        n14299), .ZN(n14292) );
  AOI222_X1 U13912 ( .A1(n16802), .A2(n13411), .B1(n16796), .B2(n13219), .C1(
        n16790), .C2(n13091), .ZN(n14299) );
  OAI221_X1 U13913 ( .B1(n7672), .B2(n16814), .C1(n7799), .C2(n16808), .A(
        n14281), .ZN(n14274) );
  AOI222_X1 U13914 ( .A1(n16802), .A2(n13410), .B1(n16796), .B2(n13218), .C1(
        n16790), .C2(n13090), .ZN(n14281) );
  OAI221_X1 U13915 ( .B1(n7670), .B2(n16814), .C1(n7797), .C2(n16808), .A(
        n14263), .ZN(n14256) );
  AOI222_X1 U13916 ( .A1(n16802), .A2(n13409), .B1(n16796), .B2(n13217), .C1(
        n16790), .C2(n13089), .ZN(n14263) );
  OAI221_X1 U13917 ( .B1(n7668), .B2(n16814), .C1(n7795), .C2(n16808), .A(
        n14245), .ZN(n14238) );
  AOI222_X1 U13918 ( .A1(n16802), .A2(n13408), .B1(n16796), .B2(n13216), .C1(
        n16790), .C2(n13088), .ZN(n14245) );
  OAI221_X1 U13919 ( .B1(n7666), .B2(n16814), .C1(n7793), .C2(n16808), .A(
        n14227), .ZN(n14220) );
  AOI222_X1 U13920 ( .A1(n16802), .A2(n13407), .B1(n16796), .B2(n13215), .C1(
        n16790), .C2(n13087), .ZN(n14227) );
  OAI221_X1 U13921 ( .B1(n7664), .B2(n16815), .C1(n7791), .C2(n16809), .A(
        n14209), .ZN(n14202) );
  AOI222_X1 U13922 ( .A1(n16803), .A2(n13406), .B1(n16797), .B2(n13214), .C1(
        n16791), .C2(n13086), .ZN(n14209) );
  OAI221_X1 U13923 ( .B1(n7662), .B2(n16815), .C1(n7789), .C2(n16809), .A(
        n14191), .ZN(n14184) );
  AOI222_X1 U13924 ( .A1(n16803), .A2(n13405), .B1(n16797), .B2(n13213), .C1(
        n16791), .C2(n13085), .ZN(n14191) );
  OAI221_X1 U13925 ( .B1(n7660), .B2(n16815), .C1(n7787), .C2(n16809), .A(
        n14173), .ZN(n14166) );
  AOI222_X1 U13926 ( .A1(n16803), .A2(n13404), .B1(n16797), .B2(n13212), .C1(
        n16791), .C2(n13084), .ZN(n14173) );
  OAI221_X1 U13927 ( .B1(n7658), .B2(n16815), .C1(n7785), .C2(n16809), .A(
        n14155), .ZN(n14148) );
  AOI222_X1 U13928 ( .A1(n16803), .A2(n13403), .B1(n16797), .B2(n13211), .C1(
        n16791), .C2(n13083), .ZN(n14155) );
  OAI221_X1 U13929 ( .B1(n7656), .B2(n16815), .C1(n7783), .C2(n16809), .A(
        n14137), .ZN(n14130) );
  AOI222_X1 U13930 ( .A1(n16803), .A2(n13402), .B1(n16797), .B2(n13210), .C1(
        n16791), .C2(n13082), .ZN(n14137) );
  OAI221_X1 U13931 ( .B1(n7654), .B2(n16815), .C1(n7781), .C2(n16809), .A(
        n14119), .ZN(n14112) );
  AOI222_X1 U13932 ( .A1(n16803), .A2(n13401), .B1(n16797), .B2(n13209), .C1(
        n16791), .C2(n13081), .ZN(n14119) );
  OAI221_X1 U13933 ( .B1(n7652), .B2(n16815), .C1(n7779), .C2(n16809), .A(
        n14101), .ZN(n14094) );
  AOI222_X1 U13934 ( .A1(n16803), .A2(n13400), .B1(n16797), .B2(n13208), .C1(
        n16791), .C2(n13080), .ZN(n14101) );
  OAI221_X1 U13935 ( .B1(n7650), .B2(n16815), .C1(n7777), .C2(n16809), .A(
        n14083), .ZN(n14076) );
  AOI222_X1 U13936 ( .A1(n16803), .A2(n13399), .B1(n16797), .B2(n13207), .C1(
        n16791), .C2(n13079), .ZN(n14083) );
  OAI221_X1 U13937 ( .B1(n7648), .B2(n16815), .C1(n7775), .C2(n16809), .A(
        n14065), .ZN(n14058) );
  AOI222_X1 U13938 ( .A1(n16803), .A2(n13398), .B1(n16797), .B2(n13206), .C1(
        n16791), .C2(n13078), .ZN(n14065) );
  OAI221_X1 U13939 ( .B1(n7646), .B2(n16815), .C1(n7773), .C2(n16809), .A(
        n14047), .ZN(n14040) );
  AOI222_X1 U13940 ( .A1(n16803), .A2(n13397), .B1(n16797), .B2(n13205), .C1(
        n16791), .C2(n13077), .ZN(n14047) );
  OAI221_X1 U13941 ( .B1(n7644), .B2(n16815), .C1(n7771), .C2(n16809), .A(
        n14029), .ZN(n14022) );
  AOI222_X1 U13942 ( .A1(n16803), .A2(n13396), .B1(n16797), .B2(n13204), .C1(
        n16791), .C2(n13076), .ZN(n14029) );
  OAI221_X1 U13943 ( .B1(n7642), .B2(n16815), .C1(n7769), .C2(n16809), .A(
        n14011), .ZN(n14004) );
  AOI222_X1 U13944 ( .A1(n16803), .A2(n13395), .B1(n16797), .B2(n13203), .C1(
        n16791), .C2(n13075), .ZN(n14011) );
  OAI221_X1 U13945 ( .B1(n7640), .B2(n16816), .C1(n7767), .C2(n16810), .A(
        n13993), .ZN(n13986) );
  AOI222_X1 U13946 ( .A1(n16804), .A2(n13394), .B1(n16798), .B2(n13202), .C1(
        n16792), .C2(n13074), .ZN(n13993) );
  OAI221_X1 U13947 ( .B1(n7638), .B2(n16816), .C1(n7765), .C2(n16810), .A(
        n13975), .ZN(n13968) );
  AOI222_X1 U13948 ( .A1(n16804), .A2(n13393), .B1(n16798), .B2(n13201), .C1(
        n16792), .C2(n13073), .ZN(n13975) );
  OAI221_X1 U13949 ( .B1(n7636), .B2(n16816), .C1(n7763), .C2(n16810), .A(
        n13957), .ZN(n13950) );
  AOI222_X1 U13950 ( .A1(n16804), .A2(n13392), .B1(n16798), .B2(n13200), .C1(
        n16792), .C2(n13072), .ZN(n13957) );
  OAI221_X1 U13951 ( .B1(n7634), .B2(n16816), .C1(n7761), .C2(n16810), .A(
        n13939), .ZN(n13932) );
  AOI222_X1 U13952 ( .A1(n16804), .A2(n13391), .B1(n16798), .B2(n13199), .C1(
        n16792), .C2(n13071), .ZN(n13939) );
  OAI221_X1 U13953 ( .B1(n7632), .B2(n16816), .C1(n7759), .C2(n16810), .A(
        n13921), .ZN(n13914) );
  AOI222_X1 U13954 ( .A1(n16804), .A2(n13390), .B1(n16798), .B2(n13198), .C1(
        n16792), .C2(n13070), .ZN(n13921) );
  OAI221_X1 U13955 ( .B1(n7630), .B2(n16816), .C1(n7757), .C2(n16810), .A(
        n13903), .ZN(n13896) );
  AOI222_X1 U13956 ( .A1(n16804), .A2(n13389), .B1(n16798), .B2(n13197), .C1(
        n16792), .C2(n13069), .ZN(n13903) );
  OAI221_X1 U13957 ( .B1(n7628), .B2(n16816), .C1(n7755), .C2(n16810), .A(
        n13885), .ZN(n13878) );
  AOI222_X1 U13958 ( .A1(n16804), .A2(n13388), .B1(n16798), .B2(n13196), .C1(
        n16792), .C2(n13068), .ZN(n13885) );
  OAI221_X1 U13959 ( .B1(n7626), .B2(n16816), .C1(n7753), .C2(n16810), .A(
        n13867), .ZN(n13860) );
  AOI222_X1 U13960 ( .A1(n16804), .A2(n13387), .B1(n16798), .B2(n13195), .C1(
        n16792), .C2(n13067), .ZN(n13867) );
  OAI221_X1 U13961 ( .B1(n7624), .B2(n16816), .C1(n7751), .C2(n16810), .A(
        n13849), .ZN(n13842) );
  AOI222_X1 U13962 ( .A1(n16804), .A2(n13386), .B1(n16798), .B2(n13194), .C1(
        n16792), .C2(n13066), .ZN(n13849) );
  OAI221_X1 U13963 ( .B1(n7622), .B2(n16816), .C1(n7749), .C2(n16810), .A(
        n13831), .ZN(n13824) );
  AOI222_X1 U13964 ( .A1(n16804), .A2(n13385), .B1(n16798), .B2(n13193), .C1(
        n16792), .C2(n13065), .ZN(n13831) );
  OAI221_X1 U13965 ( .B1(n7620), .B2(n16816), .C1(n7747), .C2(n16810), .A(
        n13813), .ZN(n13806) );
  AOI222_X1 U13966 ( .A1(n16804), .A2(n13384), .B1(n16798), .B2(n13192), .C1(
        n16792), .C2(n13064), .ZN(n13813) );
  OAI221_X1 U13967 ( .B1(n7618), .B2(n16816), .C1(n7745), .C2(n16810), .A(
        n13795), .ZN(n13788) );
  AOI222_X1 U13968 ( .A1(n16804), .A2(n13383), .B1(n16798), .B2(n13191), .C1(
        n16792), .C2(n13063), .ZN(n13795) );
  OAI221_X1 U13969 ( .B1(n13058), .B2(n16506), .C1(n964), .C2(n16500), .A(
        n16088), .ZN(n16077) );
  AOI222_X1 U13970 ( .A1(n16494), .A2(n8952), .B1(n16488), .B2(n8824), .C1(
        n16482), .C2(n8888), .ZN(n16088) );
  OAI221_X1 U13971 ( .B1(n13057), .B2(n16506), .C1(n963), .C2(n16500), .A(
        n16055), .ZN(n16048) );
  AOI222_X1 U13972 ( .A1(n16494), .A2(n8951), .B1(n16488), .B2(n8823), .C1(
        n16482), .C2(n8887), .ZN(n16055) );
  OAI221_X1 U13973 ( .B1(n13056), .B2(n16506), .C1(n962), .C2(n16500), .A(
        n16037), .ZN(n16030) );
  AOI222_X1 U13974 ( .A1(n16494), .A2(n8950), .B1(n16488), .B2(n8822), .C1(
        n16482), .C2(n8886), .ZN(n16037) );
  OAI221_X1 U13975 ( .B1(n13055), .B2(n16506), .C1(n961), .C2(n16500), .A(
        n16019), .ZN(n16012) );
  AOI222_X1 U13976 ( .A1(n16494), .A2(n8949), .B1(n16488), .B2(n8821), .C1(
        n16482), .C2(n8885), .ZN(n16019) );
  OAI221_X1 U13977 ( .B1(n13054), .B2(n16506), .C1(n960), .C2(n16500), .A(
        n16001), .ZN(n15994) );
  AOI222_X1 U13978 ( .A1(n16494), .A2(n8948), .B1(n16488), .B2(n8820), .C1(
        n16482), .C2(n8884), .ZN(n16001) );
  OAI221_X1 U13979 ( .B1(n13053), .B2(n16506), .C1(n959), .C2(n16500), .A(
        n15983), .ZN(n15976) );
  AOI222_X1 U13980 ( .A1(n16494), .A2(n8947), .B1(n16488), .B2(n8819), .C1(
        n16482), .C2(n8883), .ZN(n15983) );
  OAI221_X1 U13981 ( .B1(n13052), .B2(n16506), .C1(n958), .C2(n16500), .A(
        n15965), .ZN(n15958) );
  AOI222_X1 U13982 ( .A1(n16494), .A2(n8946), .B1(n16488), .B2(n8818), .C1(
        n16482), .C2(n8882), .ZN(n15965) );
  OAI221_X1 U13983 ( .B1(n13051), .B2(n16506), .C1(n957), .C2(n16500), .A(
        n15947), .ZN(n15940) );
  AOI222_X1 U13984 ( .A1(n16494), .A2(n8945), .B1(n16488), .B2(n8817), .C1(
        n16482), .C2(n8881), .ZN(n15947) );
  OAI221_X1 U13985 ( .B1(n13050), .B2(n16506), .C1(n956), .C2(n16500), .A(
        n15929), .ZN(n15922) );
  AOI222_X1 U13986 ( .A1(n16494), .A2(n8944), .B1(n16488), .B2(n8816), .C1(
        n16482), .C2(n8880), .ZN(n15929) );
  OAI221_X1 U13987 ( .B1(n13049), .B2(n16506), .C1(n955), .C2(n16500), .A(
        n15911), .ZN(n15904) );
  AOI222_X1 U13988 ( .A1(n16494), .A2(n8943), .B1(n16488), .B2(n8815), .C1(
        n16482), .C2(n8879), .ZN(n15911) );
  OAI221_X1 U13989 ( .B1(n13048), .B2(n16506), .C1(n954), .C2(n16500), .A(
        n15893), .ZN(n15886) );
  AOI222_X1 U13990 ( .A1(n16494), .A2(n8942), .B1(n16488), .B2(n8814), .C1(
        n16482), .C2(n8878), .ZN(n15893) );
  OAI221_X1 U13991 ( .B1(n13047), .B2(n16506), .C1(n953), .C2(n16500), .A(
        n15875), .ZN(n15868) );
  AOI222_X1 U13992 ( .A1(n16494), .A2(n8941), .B1(n16488), .B2(n8813), .C1(
        n16482), .C2(n8877), .ZN(n15875) );
  OAI221_X1 U13993 ( .B1(n13046), .B2(n16507), .C1(n952), .C2(n16501), .A(
        n15857), .ZN(n15850) );
  AOI222_X1 U13994 ( .A1(n16495), .A2(n8940), .B1(n16489), .B2(n8812), .C1(
        n16483), .C2(n8876), .ZN(n15857) );
  OAI221_X1 U13995 ( .B1(n13045), .B2(n16507), .C1(n951), .C2(n16501), .A(
        n15839), .ZN(n15832) );
  AOI222_X1 U13996 ( .A1(n16495), .A2(n8939), .B1(n16489), .B2(n8811), .C1(
        n16483), .C2(n8875), .ZN(n15839) );
  OAI221_X1 U13997 ( .B1(n13044), .B2(n16507), .C1(n950), .C2(n16501), .A(
        n15821), .ZN(n15814) );
  AOI222_X1 U13998 ( .A1(n16495), .A2(n8938), .B1(n16489), .B2(n8810), .C1(
        n16483), .C2(n8874), .ZN(n15821) );
  OAI221_X1 U13999 ( .B1(n13043), .B2(n16507), .C1(n949), .C2(n16501), .A(
        n15803), .ZN(n15796) );
  AOI222_X1 U14000 ( .A1(n16495), .A2(n8937), .B1(n16489), .B2(n8809), .C1(
        n16483), .C2(n8873), .ZN(n15803) );
  OAI221_X1 U14001 ( .B1(n13042), .B2(n16507), .C1(n948), .C2(n16501), .A(
        n15785), .ZN(n15778) );
  AOI222_X1 U14002 ( .A1(n16495), .A2(n8936), .B1(n16489), .B2(n8808), .C1(
        n16483), .C2(n8872), .ZN(n15785) );
  OAI221_X1 U14003 ( .B1(n13041), .B2(n16507), .C1(n947), .C2(n16501), .A(
        n15767), .ZN(n15760) );
  AOI222_X1 U14004 ( .A1(n16495), .A2(n8935), .B1(n16489), .B2(n8807), .C1(
        n16483), .C2(n8871), .ZN(n15767) );
  OAI221_X1 U14005 ( .B1(n13040), .B2(n16507), .C1(n946), .C2(n16501), .A(
        n15749), .ZN(n15742) );
  AOI222_X1 U14006 ( .A1(n16495), .A2(n8934), .B1(n16489), .B2(n8806), .C1(
        n16483), .C2(n8870), .ZN(n15749) );
  OAI221_X1 U14007 ( .B1(n13039), .B2(n16507), .C1(n945), .C2(n16501), .A(
        n15731), .ZN(n15724) );
  AOI222_X1 U14008 ( .A1(n16495), .A2(n8933), .B1(n16489), .B2(n8805), .C1(
        n16483), .C2(n8869), .ZN(n15731) );
  OAI221_X1 U14009 ( .B1(n13038), .B2(n16507), .C1(n944), .C2(n16501), .A(
        n15713), .ZN(n15706) );
  AOI222_X1 U14010 ( .A1(n16495), .A2(n8932), .B1(n16489), .B2(n8804), .C1(
        n16483), .C2(n8868), .ZN(n15713) );
  OAI221_X1 U14011 ( .B1(n13037), .B2(n16507), .C1(n943), .C2(n16501), .A(
        n15695), .ZN(n15688) );
  AOI222_X1 U14012 ( .A1(n16495), .A2(n8931), .B1(n16489), .B2(n8803), .C1(
        n16483), .C2(n8867), .ZN(n15695) );
  OAI221_X1 U14013 ( .B1(n13036), .B2(n16507), .C1(n942), .C2(n16501), .A(
        n15677), .ZN(n15670) );
  AOI222_X1 U14014 ( .A1(n16495), .A2(n8930), .B1(n16489), .B2(n8802), .C1(
        n16483), .C2(n8866), .ZN(n15677) );
  OAI221_X1 U14015 ( .B1(n13035), .B2(n16507), .C1(n941), .C2(n16501), .A(
        n15659), .ZN(n15652) );
  AOI222_X1 U14016 ( .A1(n16495), .A2(n8929), .B1(n16489), .B2(n8801), .C1(
        n16483), .C2(n8865), .ZN(n15659) );
  OAI221_X1 U14017 ( .B1(n13034), .B2(n16508), .C1(n940), .C2(n16502), .A(
        n15641), .ZN(n15634) );
  AOI222_X1 U14018 ( .A1(n16496), .A2(n8928), .B1(n16490), .B2(n8800), .C1(
        n16484), .C2(n8864), .ZN(n15641) );
  OAI221_X1 U14019 ( .B1(n13033), .B2(n16508), .C1(n939), .C2(n16502), .A(
        n15623), .ZN(n15616) );
  AOI222_X1 U14020 ( .A1(n16496), .A2(n8927), .B1(n16490), .B2(n8799), .C1(
        n16484), .C2(n8863), .ZN(n15623) );
  OAI221_X1 U14021 ( .B1(n13032), .B2(n16508), .C1(n938), .C2(n16502), .A(
        n15605), .ZN(n15598) );
  AOI222_X1 U14022 ( .A1(n16496), .A2(n8926), .B1(n16490), .B2(n8798), .C1(
        n16484), .C2(n8862), .ZN(n15605) );
  OAI221_X1 U14023 ( .B1(n13031), .B2(n16508), .C1(n937), .C2(n16502), .A(
        n15587), .ZN(n15580) );
  AOI222_X1 U14024 ( .A1(n16496), .A2(n8925), .B1(n16490), .B2(n8797), .C1(
        n16484), .C2(n8861), .ZN(n15587) );
  OAI221_X1 U14025 ( .B1(n13030), .B2(n16508), .C1(n936), .C2(n16502), .A(
        n15569), .ZN(n15562) );
  AOI222_X1 U14026 ( .A1(n16496), .A2(n8924), .B1(n16490), .B2(n8796), .C1(
        n16484), .C2(n8860), .ZN(n15569) );
  OAI221_X1 U14027 ( .B1(n13029), .B2(n16508), .C1(n935), .C2(n16502), .A(
        n15551), .ZN(n15544) );
  AOI222_X1 U14028 ( .A1(n16496), .A2(n8923), .B1(n16490), .B2(n8795), .C1(
        n16484), .C2(n8859), .ZN(n15551) );
  OAI221_X1 U14029 ( .B1(n13028), .B2(n16508), .C1(n934), .C2(n16502), .A(
        n15533), .ZN(n15526) );
  AOI222_X1 U14030 ( .A1(n16496), .A2(n8922), .B1(n16490), .B2(n8794), .C1(
        n16484), .C2(n8858), .ZN(n15533) );
  OAI221_X1 U14031 ( .B1(n13027), .B2(n16508), .C1(n933), .C2(n16502), .A(
        n15515), .ZN(n15508) );
  AOI222_X1 U14032 ( .A1(n16496), .A2(n8921), .B1(n16490), .B2(n8793), .C1(
        n16484), .C2(n8857), .ZN(n15515) );
  OAI221_X1 U14033 ( .B1(n13026), .B2(n16508), .C1(n932), .C2(n16502), .A(
        n15497), .ZN(n15490) );
  AOI222_X1 U14034 ( .A1(n16496), .A2(n8920), .B1(n16490), .B2(n8792), .C1(
        n16484), .C2(n8856), .ZN(n15497) );
  OAI221_X1 U14035 ( .B1(n13025), .B2(n16508), .C1(n931), .C2(n16502), .A(
        n15479), .ZN(n15472) );
  AOI222_X1 U14036 ( .A1(n16496), .A2(n8919), .B1(n16490), .B2(n8791), .C1(
        n16484), .C2(n8855), .ZN(n15479) );
  OAI221_X1 U14037 ( .B1(n13024), .B2(n16508), .C1(n930), .C2(n16502), .A(
        n15461), .ZN(n15454) );
  AOI222_X1 U14038 ( .A1(n16496), .A2(n8918), .B1(n16490), .B2(n8790), .C1(
        n16484), .C2(n8854), .ZN(n15461) );
  OAI221_X1 U14039 ( .B1(n13023), .B2(n16508), .C1(n929), .C2(n16502), .A(
        n15443), .ZN(n15436) );
  AOI222_X1 U14040 ( .A1(n16496), .A2(n8917), .B1(n16490), .B2(n8789), .C1(
        n16484), .C2(n8853), .ZN(n15443) );
  OAI221_X1 U14041 ( .B1(n13022), .B2(n16509), .C1(n928), .C2(n16503), .A(
        n15425), .ZN(n15418) );
  AOI222_X1 U14042 ( .A1(n16497), .A2(n8916), .B1(n16491), .B2(n8788), .C1(
        n16485), .C2(n8852), .ZN(n15425) );
  OAI221_X1 U14043 ( .B1(n13021), .B2(n16509), .C1(n927), .C2(n16503), .A(
        n15407), .ZN(n15400) );
  AOI222_X1 U14044 ( .A1(n16497), .A2(n8915), .B1(n16491), .B2(n8787), .C1(
        n16485), .C2(n8851), .ZN(n15407) );
  OAI221_X1 U14045 ( .B1(n13020), .B2(n16509), .C1(n926), .C2(n16503), .A(
        n15389), .ZN(n15382) );
  AOI222_X1 U14046 ( .A1(n16497), .A2(n8914), .B1(n16491), .B2(n8786), .C1(
        n16485), .C2(n8850), .ZN(n15389) );
  OAI221_X1 U14047 ( .B1(n13019), .B2(n16509), .C1(n925), .C2(n16503), .A(
        n15371), .ZN(n15364) );
  AOI222_X1 U14048 ( .A1(n16497), .A2(n8913), .B1(n16491), .B2(n8785), .C1(
        n16485), .C2(n8849), .ZN(n15371) );
  OAI221_X1 U14049 ( .B1(n13018), .B2(n16509), .C1(n924), .C2(n16503), .A(
        n15353), .ZN(n15346) );
  AOI222_X1 U14050 ( .A1(n16497), .A2(n8912), .B1(n16491), .B2(n8784), .C1(
        n16485), .C2(n8848), .ZN(n15353) );
  OAI221_X1 U14051 ( .B1(n13017), .B2(n16509), .C1(n923), .C2(n16503), .A(
        n15335), .ZN(n15328) );
  AOI222_X1 U14052 ( .A1(n16497), .A2(n8911), .B1(n16491), .B2(n8783), .C1(
        n16485), .C2(n8847), .ZN(n15335) );
  OAI221_X1 U14053 ( .B1(n13016), .B2(n16509), .C1(n922), .C2(n16503), .A(
        n15317), .ZN(n15310) );
  AOI222_X1 U14054 ( .A1(n16497), .A2(n8910), .B1(n16491), .B2(n8782), .C1(
        n16485), .C2(n8846), .ZN(n15317) );
  OAI221_X1 U14055 ( .B1(n13015), .B2(n16509), .C1(n921), .C2(n16503), .A(
        n15299), .ZN(n15292) );
  AOI222_X1 U14056 ( .A1(n16497), .A2(n8909), .B1(n16491), .B2(n8781), .C1(
        n16485), .C2(n8845), .ZN(n15299) );
  OAI221_X1 U14057 ( .B1(n13014), .B2(n16509), .C1(n920), .C2(n16503), .A(
        n15281), .ZN(n15274) );
  AOI222_X1 U14058 ( .A1(n16497), .A2(n8908), .B1(n16491), .B2(n8780), .C1(
        n16485), .C2(n8844), .ZN(n15281) );
  OAI221_X1 U14059 ( .B1(n13013), .B2(n16509), .C1(n919), .C2(n16503), .A(
        n15263), .ZN(n15256) );
  AOI222_X1 U14060 ( .A1(n16497), .A2(n8907), .B1(n16491), .B2(n8779), .C1(
        n16485), .C2(n8843), .ZN(n15263) );
  OAI221_X1 U14061 ( .B1(n13012), .B2(n16509), .C1(n918), .C2(n16503), .A(
        n15245), .ZN(n15238) );
  AOI222_X1 U14062 ( .A1(n16497), .A2(n8906), .B1(n16491), .B2(n8778), .C1(
        n16485), .C2(n8842), .ZN(n15245) );
  OAI221_X1 U14063 ( .B1(n13011), .B2(n16509), .C1(n917), .C2(n16503), .A(
        n15227), .ZN(n15220) );
  AOI222_X1 U14064 ( .A1(n16497), .A2(n8905), .B1(n16491), .B2(n8777), .C1(
        n16485), .C2(n8841), .ZN(n15227) );
  OAI221_X1 U14065 ( .B1(n13058), .B2(n16711), .C1(n964), .C2(n16705), .A(
        n14880), .ZN(n14869) );
  AOI222_X1 U14066 ( .A1(n16699), .A2(n8952), .B1(n16693), .B2(n8824), .C1(
        n16687), .C2(n8888), .ZN(n14880) );
  OAI221_X1 U14067 ( .B1(n13057), .B2(n16711), .C1(n963), .C2(n16705), .A(
        n14847), .ZN(n14840) );
  AOI222_X1 U14068 ( .A1(n16699), .A2(n8951), .B1(n16693), .B2(n8823), .C1(
        n16687), .C2(n8887), .ZN(n14847) );
  OAI221_X1 U14069 ( .B1(n13056), .B2(n16711), .C1(n962), .C2(n16705), .A(
        n14829), .ZN(n14822) );
  AOI222_X1 U14070 ( .A1(n16699), .A2(n8950), .B1(n16693), .B2(n8822), .C1(
        n16687), .C2(n8886), .ZN(n14829) );
  OAI221_X1 U14071 ( .B1(n13055), .B2(n16711), .C1(n961), .C2(n16705), .A(
        n14811), .ZN(n14804) );
  AOI222_X1 U14072 ( .A1(n16699), .A2(n8949), .B1(n16693), .B2(n8821), .C1(
        n16687), .C2(n8885), .ZN(n14811) );
  OAI221_X1 U14073 ( .B1(n13054), .B2(n16711), .C1(n960), .C2(n16705), .A(
        n14793), .ZN(n14786) );
  AOI222_X1 U14074 ( .A1(n16699), .A2(n8948), .B1(n16693), .B2(n8820), .C1(
        n16687), .C2(n8884), .ZN(n14793) );
  OAI221_X1 U14075 ( .B1(n13053), .B2(n16711), .C1(n959), .C2(n16705), .A(
        n14775), .ZN(n14768) );
  AOI222_X1 U14076 ( .A1(n16699), .A2(n8947), .B1(n16693), .B2(n8819), .C1(
        n16687), .C2(n8883), .ZN(n14775) );
  OAI221_X1 U14077 ( .B1(n13052), .B2(n16711), .C1(n958), .C2(n16705), .A(
        n14757), .ZN(n14750) );
  AOI222_X1 U14078 ( .A1(n16699), .A2(n8946), .B1(n16693), .B2(n8818), .C1(
        n16687), .C2(n8882), .ZN(n14757) );
  OAI221_X1 U14079 ( .B1(n13051), .B2(n16711), .C1(n957), .C2(n16705), .A(
        n14739), .ZN(n14732) );
  AOI222_X1 U14080 ( .A1(n16699), .A2(n8945), .B1(n16693), .B2(n8817), .C1(
        n16687), .C2(n8881), .ZN(n14739) );
  OAI221_X1 U14081 ( .B1(n13050), .B2(n16711), .C1(n956), .C2(n16705), .A(
        n14721), .ZN(n14714) );
  AOI222_X1 U14082 ( .A1(n16699), .A2(n8944), .B1(n16693), .B2(n8816), .C1(
        n16687), .C2(n8880), .ZN(n14721) );
  OAI221_X1 U14083 ( .B1(n13049), .B2(n16711), .C1(n955), .C2(n16705), .A(
        n14703), .ZN(n14696) );
  AOI222_X1 U14084 ( .A1(n16699), .A2(n8943), .B1(n16693), .B2(n8815), .C1(
        n16687), .C2(n8879), .ZN(n14703) );
  OAI221_X1 U14085 ( .B1(n13048), .B2(n16711), .C1(n954), .C2(n16705), .A(
        n14685), .ZN(n14678) );
  AOI222_X1 U14086 ( .A1(n16699), .A2(n8942), .B1(n16693), .B2(n8814), .C1(
        n16687), .C2(n8878), .ZN(n14685) );
  OAI221_X1 U14087 ( .B1(n13047), .B2(n16711), .C1(n953), .C2(n16705), .A(
        n14667), .ZN(n14660) );
  AOI222_X1 U14088 ( .A1(n16699), .A2(n8941), .B1(n16693), .B2(n8813), .C1(
        n16687), .C2(n8877), .ZN(n14667) );
  OAI221_X1 U14089 ( .B1(n13046), .B2(n16712), .C1(n952), .C2(n16706), .A(
        n14649), .ZN(n14642) );
  AOI222_X1 U14090 ( .A1(n16700), .A2(n8940), .B1(n16694), .B2(n8812), .C1(
        n16688), .C2(n8876), .ZN(n14649) );
  OAI221_X1 U14091 ( .B1(n13045), .B2(n16712), .C1(n951), .C2(n16706), .A(
        n14631), .ZN(n14624) );
  AOI222_X1 U14092 ( .A1(n16700), .A2(n8939), .B1(n16694), .B2(n8811), .C1(
        n16688), .C2(n8875), .ZN(n14631) );
  OAI221_X1 U14093 ( .B1(n13044), .B2(n16712), .C1(n950), .C2(n16706), .A(
        n14613), .ZN(n14606) );
  AOI222_X1 U14094 ( .A1(n16700), .A2(n8938), .B1(n16694), .B2(n8810), .C1(
        n16688), .C2(n8874), .ZN(n14613) );
  OAI221_X1 U14095 ( .B1(n13043), .B2(n16712), .C1(n949), .C2(n16706), .A(
        n14595), .ZN(n14588) );
  AOI222_X1 U14096 ( .A1(n16700), .A2(n8937), .B1(n16694), .B2(n8809), .C1(
        n16688), .C2(n8873), .ZN(n14595) );
  OAI221_X1 U14097 ( .B1(n13042), .B2(n16712), .C1(n948), .C2(n16706), .A(
        n14577), .ZN(n14570) );
  AOI222_X1 U14098 ( .A1(n16700), .A2(n8936), .B1(n16694), .B2(n8808), .C1(
        n16688), .C2(n8872), .ZN(n14577) );
  OAI221_X1 U14099 ( .B1(n13041), .B2(n16712), .C1(n947), .C2(n16706), .A(
        n14559), .ZN(n14552) );
  AOI222_X1 U14100 ( .A1(n16700), .A2(n8935), .B1(n16694), .B2(n8807), .C1(
        n16688), .C2(n8871), .ZN(n14559) );
  OAI221_X1 U14101 ( .B1(n13040), .B2(n16712), .C1(n946), .C2(n16706), .A(
        n14541), .ZN(n14534) );
  AOI222_X1 U14102 ( .A1(n16700), .A2(n8934), .B1(n16694), .B2(n8806), .C1(
        n16688), .C2(n8870), .ZN(n14541) );
  OAI221_X1 U14103 ( .B1(n13039), .B2(n16712), .C1(n945), .C2(n16706), .A(
        n14523), .ZN(n14516) );
  AOI222_X1 U14104 ( .A1(n16700), .A2(n8933), .B1(n16694), .B2(n8805), .C1(
        n16688), .C2(n8869), .ZN(n14523) );
  OAI221_X1 U14105 ( .B1(n13038), .B2(n16712), .C1(n944), .C2(n16706), .A(
        n14505), .ZN(n14498) );
  AOI222_X1 U14106 ( .A1(n16700), .A2(n8932), .B1(n16694), .B2(n8804), .C1(
        n16688), .C2(n8868), .ZN(n14505) );
  OAI221_X1 U14107 ( .B1(n13037), .B2(n16712), .C1(n943), .C2(n16706), .A(
        n14487), .ZN(n14480) );
  AOI222_X1 U14108 ( .A1(n16700), .A2(n8931), .B1(n16694), .B2(n8803), .C1(
        n16688), .C2(n8867), .ZN(n14487) );
  OAI221_X1 U14109 ( .B1(n13036), .B2(n16712), .C1(n942), .C2(n16706), .A(
        n14469), .ZN(n14462) );
  AOI222_X1 U14110 ( .A1(n16700), .A2(n8930), .B1(n16694), .B2(n8802), .C1(
        n16688), .C2(n8866), .ZN(n14469) );
  OAI221_X1 U14111 ( .B1(n13035), .B2(n16712), .C1(n941), .C2(n16706), .A(
        n14451), .ZN(n14444) );
  AOI222_X1 U14112 ( .A1(n16700), .A2(n8929), .B1(n16694), .B2(n8801), .C1(
        n16688), .C2(n8865), .ZN(n14451) );
  OAI221_X1 U14113 ( .B1(n13034), .B2(n16713), .C1(n940), .C2(n16707), .A(
        n14433), .ZN(n14426) );
  AOI222_X1 U14114 ( .A1(n16701), .A2(n8928), .B1(n16695), .B2(n8800), .C1(
        n16689), .C2(n8864), .ZN(n14433) );
  OAI221_X1 U14115 ( .B1(n13033), .B2(n16713), .C1(n939), .C2(n16707), .A(
        n14415), .ZN(n14408) );
  AOI222_X1 U14116 ( .A1(n16701), .A2(n8927), .B1(n16695), .B2(n8799), .C1(
        n16689), .C2(n8863), .ZN(n14415) );
  OAI221_X1 U14117 ( .B1(n13032), .B2(n16713), .C1(n938), .C2(n16707), .A(
        n14397), .ZN(n14390) );
  AOI222_X1 U14118 ( .A1(n16701), .A2(n8926), .B1(n16695), .B2(n8798), .C1(
        n16689), .C2(n8862), .ZN(n14397) );
  OAI221_X1 U14119 ( .B1(n13031), .B2(n16713), .C1(n937), .C2(n16707), .A(
        n14379), .ZN(n14372) );
  AOI222_X1 U14120 ( .A1(n16701), .A2(n8925), .B1(n16695), .B2(n8797), .C1(
        n16689), .C2(n8861), .ZN(n14379) );
  OAI221_X1 U14121 ( .B1(n13030), .B2(n16713), .C1(n936), .C2(n16707), .A(
        n14361), .ZN(n14354) );
  AOI222_X1 U14122 ( .A1(n16701), .A2(n8924), .B1(n16695), .B2(n8796), .C1(
        n16689), .C2(n8860), .ZN(n14361) );
  OAI221_X1 U14123 ( .B1(n13029), .B2(n16713), .C1(n935), .C2(n16707), .A(
        n14343), .ZN(n14336) );
  AOI222_X1 U14124 ( .A1(n16701), .A2(n8923), .B1(n16695), .B2(n8795), .C1(
        n16689), .C2(n8859), .ZN(n14343) );
  OAI221_X1 U14125 ( .B1(n13028), .B2(n16713), .C1(n934), .C2(n16707), .A(
        n14325), .ZN(n14318) );
  AOI222_X1 U14126 ( .A1(n16701), .A2(n8922), .B1(n16695), .B2(n8794), .C1(
        n16689), .C2(n8858), .ZN(n14325) );
  OAI221_X1 U14127 ( .B1(n13027), .B2(n16713), .C1(n933), .C2(n16707), .A(
        n14307), .ZN(n14300) );
  AOI222_X1 U14128 ( .A1(n16701), .A2(n8921), .B1(n16695), .B2(n8793), .C1(
        n16689), .C2(n8857), .ZN(n14307) );
  OAI221_X1 U14129 ( .B1(n13026), .B2(n16713), .C1(n932), .C2(n16707), .A(
        n14289), .ZN(n14282) );
  AOI222_X1 U14130 ( .A1(n16701), .A2(n8920), .B1(n16695), .B2(n8792), .C1(
        n16689), .C2(n8856), .ZN(n14289) );
  OAI221_X1 U14131 ( .B1(n13025), .B2(n16713), .C1(n931), .C2(n16707), .A(
        n14271), .ZN(n14264) );
  AOI222_X1 U14132 ( .A1(n16701), .A2(n8919), .B1(n16695), .B2(n8791), .C1(
        n16689), .C2(n8855), .ZN(n14271) );
  OAI221_X1 U14133 ( .B1(n13024), .B2(n16713), .C1(n930), .C2(n16707), .A(
        n14253), .ZN(n14246) );
  AOI222_X1 U14134 ( .A1(n16701), .A2(n8918), .B1(n16695), .B2(n8790), .C1(
        n16689), .C2(n8854), .ZN(n14253) );
  OAI221_X1 U14135 ( .B1(n13023), .B2(n16713), .C1(n929), .C2(n16707), .A(
        n14235), .ZN(n14228) );
  AOI222_X1 U14136 ( .A1(n16701), .A2(n8917), .B1(n16695), .B2(n8789), .C1(
        n16689), .C2(n8853), .ZN(n14235) );
  OAI221_X1 U14137 ( .B1(n13022), .B2(n16714), .C1(n928), .C2(n16708), .A(
        n14217), .ZN(n14210) );
  AOI222_X1 U14138 ( .A1(n16702), .A2(n8916), .B1(n16696), .B2(n8788), .C1(
        n16690), .C2(n8852), .ZN(n14217) );
  OAI221_X1 U14139 ( .B1(n13021), .B2(n16714), .C1(n927), .C2(n16708), .A(
        n14199), .ZN(n14192) );
  AOI222_X1 U14140 ( .A1(n16702), .A2(n8915), .B1(n16696), .B2(n8787), .C1(
        n16690), .C2(n8851), .ZN(n14199) );
  OAI221_X1 U14141 ( .B1(n13020), .B2(n16714), .C1(n926), .C2(n16708), .A(
        n14181), .ZN(n14174) );
  AOI222_X1 U14142 ( .A1(n16702), .A2(n8914), .B1(n16696), .B2(n8786), .C1(
        n16690), .C2(n8850), .ZN(n14181) );
  OAI221_X1 U14143 ( .B1(n13019), .B2(n16714), .C1(n925), .C2(n16708), .A(
        n14163), .ZN(n14156) );
  AOI222_X1 U14144 ( .A1(n16702), .A2(n8913), .B1(n16696), .B2(n8785), .C1(
        n16690), .C2(n8849), .ZN(n14163) );
  OAI221_X1 U14145 ( .B1(n13018), .B2(n16714), .C1(n924), .C2(n16708), .A(
        n14145), .ZN(n14138) );
  AOI222_X1 U14146 ( .A1(n16702), .A2(n8912), .B1(n16696), .B2(n8784), .C1(
        n16690), .C2(n8848), .ZN(n14145) );
  OAI221_X1 U14147 ( .B1(n13017), .B2(n16714), .C1(n923), .C2(n16708), .A(
        n14127), .ZN(n14120) );
  AOI222_X1 U14148 ( .A1(n16702), .A2(n8911), .B1(n16696), .B2(n8783), .C1(
        n16690), .C2(n8847), .ZN(n14127) );
  OAI221_X1 U14149 ( .B1(n13016), .B2(n16714), .C1(n922), .C2(n16708), .A(
        n14109), .ZN(n14102) );
  AOI222_X1 U14150 ( .A1(n16702), .A2(n8910), .B1(n16696), .B2(n8782), .C1(
        n16690), .C2(n8846), .ZN(n14109) );
  OAI221_X1 U14151 ( .B1(n13015), .B2(n16714), .C1(n921), .C2(n16708), .A(
        n14091), .ZN(n14084) );
  AOI222_X1 U14152 ( .A1(n16702), .A2(n8909), .B1(n16696), .B2(n8781), .C1(
        n16690), .C2(n8845), .ZN(n14091) );
  OAI221_X1 U14153 ( .B1(n13014), .B2(n16714), .C1(n920), .C2(n16708), .A(
        n14073), .ZN(n14066) );
  AOI222_X1 U14154 ( .A1(n16702), .A2(n8908), .B1(n16696), .B2(n8780), .C1(
        n16690), .C2(n8844), .ZN(n14073) );
  OAI221_X1 U14155 ( .B1(n13013), .B2(n16714), .C1(n919), .C2(n16708), .A(
        n14055), .ZN(n14048) );
  AOI222_X1 U14156 ( .A1(n16702), .A2(n8907), .B1(n16696), .B2(n8779), .C1(
        n16690), .C2(n8843), .ZN(n14055) );
  OAI221_X1 U14157 ( .B1(n13012), .B2(n16714), .C1(n918), .C2(n16708), .A(
        n14037), .ZN(n14030) );
  AOI222_X1 U14158 ( .A1(n16702), .A2(n8906), .B1(n16696), .B2(n8778), .C1(
        n16690), .C2(n8842), .ZN(n14037) );
  OAI221_X1 U14159 ( .B1(n13011), .B2(n16714), .C1(n917), .C2(n16708), .A(
        n14019), .ZN(n14012) );
  AOI222_X1 U14160 ( .A1(n16702), .A2(n8905), .B1(n16696), .B2(n8777), .C1(
        n16690), .C2(n8841), .ZN(n14019) );
  OAI221_X1 U14161 ( .B1(n13010), .B2(n16510), .C1(n916), .C2(n16504), .A(
        n15209), .ZN(n15202) );
  AOI222_X1 U14162 ( .A1(n16498), .A2(n8904), .B1(n16492), .B2(n8776), .C1(
        n16486), .C2(n8840), .ZN(n15209) );
  OAI221_X1 U14163 ( .B1(n13009), .B2(n16510), .C1(n915), .C2(n16504), .A(
        n15191), .ZN(n15184) );
  AOI222_X1 U14164 ( .A1(n16498), .A2(n8903), .B1(n16492), .B2(n8775), .C1(
        n16486), .C2(n8839), .ZN(n15191) );
  OAI221_X1 U14165 ( .B1(n13008), .B2(n16510), .C1(n914), .C2(n16504), .A(
        n15173), .ZN(n15166) );
  AOI222_X1 U14166 ( .A1(n16498), .A2(n8902), .B1(n16492), .B2(n8774), .C1(
        n16486), .C2(n8838), .ZN(n15173) );
  OAI221_X1 U14167 ( .B1(n13007), .B2(n16510), .C1(n913), .C2(n16504), .A(
        n15155), .ZN(n15148) );
  AOI222_X1 U14168 ( .A1(n16498), .A2(n8901), .B1(n16492), .B2(n8773), .C1(
        n16486), .C2(n8837), .ZN(n15155) );
  OAI221_X1 U14169 ( .B1(n13006), .B2(n16510), .C1(n912), .C2(n16504), .A(
        n15137), .ZN(n15130) );
  AOI222_X1 U14170 ( .A1(n16498), .A2(n8900), .B1(n16492), .B2(n8772), .C1(
        n16486), .C2(n8836), .ZN(n15137) );
  OAI221_X1 U14171 ( .B1(n13005), .B2(n16510), .C1(n911), .C2(n16504), .A(
        n15119), .ZN(n15112) );
  AOI222_X1 U14172 ( .A1(n16498), .A2(n8899), .B1(n16492), .B2(n8771), .C1(
        n16486), .C2(n8835), .ZN(n15119) );
  OAI221_X1 U14173 ( .B1(n13004), .B2(n16510), .C1(n910), .C2(n16504), .A(
        n15101), .ZN(n15094) );
  AOI222_X1 U14174 ( .A1(n16498), .A2(n8898), .B1(n16492), .B2(n8770), .C1(
        n16486), .C2(n8834), .ZN(n15101) );
  OAI221_X1 U14175 ( .B1(n13003), .B2(n16510), .C1(n909), .C2(n16504), .A(
        n15083), .ZN(n15076) );
  AOI222_X1 U14176 ( .A1(n16498), .A2(n8897), .B1(n16492), .B2(n8769), .C1(
        n16486), .C2(n8833), .ZN(n15083) );
  OAI221_X1 U14177 ( .B1(n13002), .B2(n16510), .C1(n908), .C2(n16504), .A(
        n15065), .ZN(n15058) );
  AOI222_X1 U14178 ( .A1(n16498), .A2(n8896), .B1(n16492), .B2(n8768), .C1(
        n16486), .C2(n8832), .ZN(n15065) );
  OAI221_X1 U14179 ( .B1(n13001), .B2(n16510), .C1(n907), .C2(n16504), .A(
        n15047), .ZN(n15040) );
  AOI222_X1 U14180 ( .A1(n16498), .A2(n8895), .B1(n16492), .B2(n8767), .C1(
        n16486), .C2(n8831), .ZN(n15047) );
  OAI221_X1 U14181 ( .B1(n13000), .B2(n16510), .C1(n906), .C2(n16504), .A(
        n15029), .ZN(n15022) );
  AOI222_X1 U14182 ( .A1(n16498), .A2(n8894), .B1(n16492), .B2(n8766), .C1(
        n16486), .C2(n8830), .ZN(n15029) );
  OAI221_X1 U14183 ( .B1(n12999), .B2(n16510), .C1(n905), .C2(n16504), .A(
        n15011), .ZN(n15004) );
  AOI222_X1 U14184 ( .A1(n16498), .A2(n8893), .B1(n16492), .B2(n8765), .C1(
        n16486), .C2(n8829), .ZN(n15011) );
  OAI221_X1 U14185 ( .B1(n13010), .B2(n16715), .C1(n916), .C2(n16709), .A(
        n14001), .ZN(n13994) );
  AOI222_X1 U14186 ( .A1(n16703), .A2(n8904), .B1(n16697), .B2(n8776), .C1(
        n16691), .C2(n8840), .ZN(n14001) );
  OAI221_X1 U14187 ( .B1(n13009), .B2(n16715), .C1(n915), .C2(n16709), .A(
        n13983), .ZN(n13976) );
  AOI222_X1 U14188 ( .A1(n16703), .A2(n8903), .B1(n16697), .B2(n8775), .C1(
        n16691), .C2(n8839), .ZN(n13983) );
  OAI221_X1 U14189 ( .B1(n13008), .B2(n16715), .C1(n914), .C2(n16709), .A(
        n13965), .ZN(n13958) );
  AOI222_X1 U14190 ( .A1(n16703), .A2(n8902), .B1(n16697), .B2(n8774), .C1(
        n16691), .C2(n8838), .ZN(n13965) );
  OAI221_X1 U14191 ( .B1(n13007), .B2(n16715), .C1(n913), .C2(n16709), .A(
        n13947), .ZN(n13940) );
  AOI222_X1 U14192 ( .A1(n16703), .A2(n8901), .B1(n16697), .B2(n8773), .C1(
        n16691), .C2(n8837), .ZN(n13947) );
  OAI221_X1 U14193 ( .B1(n13006), .B2(n16715), .C1(n912), .C2(n16709), .A(
        n13929), .ZN(n13922) );
  AOI222_X1 U14194 ( .A1(n16703), .A2(n8900), .B1(n16697), .B2(n8772), .C1(
        n16691), .C2(n8836), .ZN(n13929) );
  OAI221_X1 U14195 ( .B1(n13005), .B2(n16715), .C1(n911), .C2(n16709), .A(
        n13911), .ZN(n13904) );
  AOI222_X1 U14196 ( .A1(n16703), .A2(n8899), .B1(n16697), .B2(n8771), .C1(
        n16691), .C2(n8835), .ZN(n13911) );
  OAI221_X1 U14197 ( .B1(n13004), .B2(n16715), .C1(n910), .C2(n16709), .A(
        n13893), .ZN(n13886) );
  AOI222_X1 U14198 ( .A1(n16703), .A2(n8898), .B1(n16697), .B2(n8770), .C1(
        n16691), .C2(n8834), .ZN(n13893) );
  OAI221_X1 U14199 ( .B1(n13003), .B2(n16715), .C1(n909), .C2(n16709), .A(
        n13875), .ZN(n13868) );
  AOI222_X1 U14200 ( .A1(n16703), .A2(n8897), .B1(n16697), .B2(n8769), .C1(
        n16691), .C2(n8833), .ZN(n13875) );
  OAI221_X1 U14201 ( .B1(n13002), .B2(n16715), .C1(n908), .C2(n16709), .A(
        n13857), .ZN(n13850) );
  AOI222_X1 U14202 ( .A1(n16703), .A2(n8896), .B1(n16697), .B2(n8768), .C1(
        n16691), .C2(n8832), .ZN(n13857) );
  OAI221_X1 U14203 ( .B1(n13001), .B2(n16715), .C1(n907), .C2(n16709), .A(
        n13839), .ZN(n13832) );
  AOI222_X1 U14204 ( .A1(n16703), .A2(n8895), .B1(n16697), .B2(n8767), .C1(
        n16691), .C2(n8831), .ZN(n13839) );
  OAI221_X1 U14205 ( .B1(n13000), .B2(n16715), .C1(n906), .C2(n16709), .A(
        n13821), .ZN(n13814) );
  AOI222_X1 U14206 ( .A1(n16703), .A2(n8894), .B1(n16697), .B2(n8766), .C1(
        n16691), .C2(n8830), .ZN(n13821) );
  OAI221_X1 U14207 ( .B1(n12999), .B2(n16715), .C1(n905), .C2(n16709), .A(
        n13803), .ZN(n13796) );
  AOI222_X1 U14208 ( .A1(n16703), .A2(n8893), .B1(n16697), .B2(n8765), .C1(
        n16691), .C2(n8829), .ZN(n13803) );
  OAI22_X1 U14209 ( .A1(n16961), .A2(n17432), .B1(n16959), .B2(n13378), .ZN(
        n5260) );
  OAI22_X1 U14210 ( .A1(n16961), .A2(n17434), .B1(n16959), .B2(n13377), .ZN(
        n5261) );
  OAI22_X1 U14211 ( .A1(n16961), .A2(n17436), .B1(n16959), .B2(n13376), .ZN(
        n5262) );
  OAI22_X1 U14212 ( .A1(n16961), .A2(n17438), .B1(n16959), .B2(n13375), .ZN(
        n5263) );
  OAI22_X1 U14213 ( .A1(n16961), .A2(n17440), .B1(n16959), .B2(n13374), .ZN(
        n5264) );
  OAI22_X1 U14214 ( .A1(n16962), .A2(n17442), .B1(n16959), .B2(n13373), .ZN(
        n5265) );
  OAI22_X1 U14215 ( .A1(n16962), .A2(n17444), .B1(n16959), .B2(n13372), .ZN(
        n5266) );
  OAI22_X1 U14216 ( .A1(n16962), .A2(n17446), .B1(n16959), .B2(n13371), .ZN(
        n5267) );
  OAI22_X1 U14217 ( .A1(n16962), .A2(n17448), .B1(n16959), .B2(n13370), .ZN(
        n5268) );
  OAI22_X1 U14218 ( .A1(n16962), .A2(n17450), .B1(n16959), .B2(n13369), .ZN(
        n5269) );
  OAI22_X1 U14219 ( .A1(n16963), .A2(n17452), .B1(n16959), .B2(n13368), .ZN(
        n5270) );
  OAI22_X1 U14220 ( .A1(n16963), .A2(n17454), .B1(n16959), .B2(n13367), .ZN(
        n5271) );
  OAI22_X1 U14221 ( .A1(n16963), .A2(n17456), .B1(n16960), .B2(n13366), .ZN(
        n5272) );
  OAI22_X1 U14222 ( .A1(n16963), .A2(n17458), .B1(n16960), .B2(n13365), .ZN(
        n5273) );
  OAI22_X1 U14223 ( .A1(n16963), .A2(n17460), .B1(n16960), .B2(n13364), .ZN(
        n5274) );
  OAI22_X1 U14224 ( .A1(n16964), .A2(n17462), .B1(n16960), .B2(n13363), .ZN(
        n5275) );
  OAI22_X1 U14225 ( .A1(n16964), .A2(n17464), .B1(n16960), .B2(n13362), .ZN(
        n5276) );
  OAI22_X1 U14226 ( .A1(n16964), .A2(n17466), .B1(n16960), .B2(n13361), .ZN(
        n5277) );
  OAI22_X1 U14227 ( .A1(n16964), .A2(n17468), .B1(n16960), .B2(n13360), .ZN(
        n5278) );
  OAI22_X1 U14228 ( .A1(n16964), .A2(n17470), .B1(n16960), .B2(n13359), .ZN(
        n5279) );
  OAI22_X1 U14229 ( .A1(n16965), .A2(n17472), .B1(n16960), .B2(n13358), .ZN(
        n5280) );
  OAI22_X1 U14230 ( .A1(n16965), .A2(n17474), .B1(n16960), .B2(n13357), .ZN(
        n5281) );
  OAI22_X1 U14231 ( .A1(n16965), .A2(n17476), .B1(n16960), .B2(n13356), .ZN(
        n5282) );
  OAI22_X1 U14232 ( .A1(n16965), .A2(n17478), .B1(n16960), .B2(n13355), .ZN(
        n5283) );
  OAI22_X1 U14233 ( .A1(n16978), .A2(n17432), .B1(n16976), .B2(n13314), .ZN(
        n5324) );
  OAI22_X1 U14234 ( .A1(n16978), .A2(n17434), .B1(n16976), .B2(n13313), .ZN(
        n5325) );
  OAI22_X1 U14235 ( .A1(n16978), .A2(n17436), .B1(n16976), .B2(n13312), .ZN(
        n5326) );
  OAI22_X1 U14236 ( .A1(n16978), .A2(n17438), .B1(n16976), .B2(n13311), .ZN(
        n5327) );
  OAI22_X1 U14237 ( .A1(n16978), .A2(n17440), .B1(n16976), .B2(n13310), .ZN(
        n5328) );
  OAI22_X1 U14238 ( .A1(n16979), .A2(n17442), .B1(n16976), .B2(n13309), .ZN(
        n5329) );
  OAI22_X1 U14239 ( .A1(n16979), .A2(n17444), .B1(n16976), .B2(n13308), .ZN(
        n5330) );
  OAI22_X1 U14240 ( .A1(n16979), .A2(n17446), .B1(n16976), .B2(n13307), .ZN(
        n5331) );
  OAI22_X1 U14241 ( .A1(n16979), .A2(n17448), .B1(n16976), .B2(n13306), .ZN(
        n5332) );
  OAI22_X1 U14242 ( .A1(n16979), .A2(n17450), .B1(n16976), .B2(n13305), .ZN(
        n5333) );
  OAI22_X1 U14243 ( .A1(n16980), .A2(n17452), .B1(n16976), .B2(n13304), .ZN(
        n5334) );
  OAI22_X1 U14244 ( .A1(n16980), .A2(n17454), .B1(n16976), .B2(n13303), .ZN(
        n5335) );
  OAI22_X1 U14245 ( .A1(n16980), .A2(n17456), .B1(n16977), .B2(n13302), .ZN(
        n5336) );
  OAI22_X1 U14246 ( .A1(n16980), .A2(n17458), .B1(n16977), .B2(n13301), .ZN(
        n5337) );
  OAI22_X1 U14247 ( .A1(n16980), .A2(n17460), .B1(n16977), .B2(n13300), .ZN(
        n5338) );
  OAI22_X1 U14248 ( .A1(n16981), .A2(n17462), .B1(n16977), .B2(n13299), .ZN(
        n5339) );
  OAI22_X1 U14249 ( .A1(n16981), .A2(n17464), .B1(n16977), .B2(n13298), .ZN(
        n5340) );
  OAI22_X1 U14250 ( .A1(n16981), .A2(n17466), .B1(n16977), .B2(n13297), .ZN(
        n5341) );
  OAI22_X1 U14251 ( .A1(n16981), .A2(n17468), .B1(n16977), .B2(n13296), .ZN(
        n5342) );
  OAI22_X1 U14252 ( .A1(n16981), .A2(n17470), .B1(n16977), .B2(n13295), .ZN(
        n5343) );
  OAI22_X1 U14253 ( .A1(n16982), .A2(n17472), .B1(n16977), .B2(n13294), .ZN(
        n5344) );
  OAI22_X1 U14254 ( .A1(n16982), .A2(n17474), .B1(n16977), .B2(n13293), .ZN(
        n5345) );
  OAI22_X1 U14255 ( .A1(n16982), .A2(n17476), .B1(n16977), .B2(n13292), .ZN(
        n5346) );
  OAI22_X1 U14256 ( .A1(n16982), .A2(n17478), .B1(n16977), .B2(n13291), .ZN(
        n5347) );
  OAI22_X1 U14257 ( .A1(n17080), .A2(n17432), .B1(n17078), .B2(n12994), .ZN(
        n5708) );
  OAI22_X1 U14258 ( .A1(n17080), .A2(n17434), .B1(n17078), .B2(n12993), .ZN(
        n5709) );
  OAI22_X1 U14259 ( .A1(n17080), .A2(n17436), .B1(n17078), .B2(n12992), .ZN(
        n5710) );
  OAI22_X1 U14260 ( .A1(n17080), .A2(n17438), .B1(n17078), .B2(n12991), .ZN(
        n5711) );
  OAI22_X1 U14261 ( .A1(n17080), .A2(n17440), .B1(n17078), .B2(n12990), .ZN(
        n5712) );
  OAI22_X1 U14262 ( .A1(n17081), .A2(n17442), .B1(n17078), .B2(n12989), .ZN(
        n5713) );
  OAI22_X1 U14263 ( .A1(n17081), .A2(n17444), .B1(n17078), .B2(n12988), .ZN(
        n5714) );
  OAI22_X1 U14264 ( .A1(n17081), .A2(n17446), .B1(n17078), .B2(n12987), .ZN(
        n5715) );
  OAI22_X1 U14265 ( .A1(n17081), .A2(n17448), .B1(n17078), .B2(n12986), .ZN(
        n5716) );
  OAI22_X1 U14266 ( .A1(n17081), .A2(n17450), .B1(n17078), .B2(n12985), .ZN(
        n5717) );
  OAI22_X1 U14267 ( .A1(n17082), .A2(n17452), .B1(n17078), .B2(n12984), .ZN(
        n5718) );
  OAI22_X1 U14268 ( .A1(n17082), .A2(n17454), .B1(n17078), .B2(n12983), .ZN(
        n5719) );
  OAI22_X1 U14269 ( .A1(n17082), .A2(n17456), .B1(n17079), .B2(n12982), .ZN(
        n5720) );
  OAI22_X1 U14270 ( .A1(n17082), .A2(n17458), .B1(n17079), .B2(n12981), .ZN(
        n5721) );
  OAI22_X1 U14271 ( .A1(n17082), .A2(n17460), .B1(n17079), .B2(n12980), .ZN(
        n5722) );
  OAI22_X1 U14272 ( .A1(n17083), .A2(n17462), .B1(n17079), .B2(n12979), .ZN(
        n5723) );
  OAI22_X1 U14273 ( .A1(n17083), .A2(n17464), .B1(n17079), .B2(n12978), .ZN(
        n5724) );
  OAI22_X1 U14274 ( .A1(n17083), .A2(n17466), .B1(n17079), .B2(n12977), .ZN(
        n5725) );
  OAI22_X1 U14275 ( .A1(n17083), .A2(n17468), .B1(n17079), .B2(n12976), .ZN(
        n5726) );
  OAI22_X1 U14276 ( .A1(n17083), .A2(n17470), .B1(n17079), .B2(n12975), .ZN(
        n5727) );
  OAI22_X1 U14277 ( .A1(n17084), .A2(n17472), .B1(n17079), .B2(n12974), .ZN(
        n5728) );
  OAI22_X1 U14278 ( .A1(n17084), .A2(n17474), .B1(n17079), .B2(n12973), .ZN(
        n5729) );
  OAI22_X1 U14279 ( .A1(n17084), .A2(n17476), .B1(n17079), .B2(n12972), .ZN(
        n5730) );
  OAI22_X1 U14280 ( .A1(n17084), .A2(n17478), .B1(n17079), .B2(n12971), .ZN(
        n5731) );
  OAI22_X1 U14281 ( .A1(n17131), .A2(n17433), .B1(n17129), .B2(n12930), .ZN(
        n5900) );
  OAI22_X1 U14282 ( .A1(n17131), .A2(n17435), .B1(n17129), .B2(n12929), .ZN(
        n5901) );
  OAI22_X1 U14283 ( .A1(n17131), .A2(n17437), .B1(n17129), .B2(n12928), .ZN(
        n5902) );
  OAI22_X1 U14284 ( .A1(n17131), .A2(n17439), .B1(n17129), .B2(n12927), .ZN(
        n5903) );
  OAI22_X1 U14285 ( .A1(n17131), .A2(n17441), .B1(n17129), .B2(n12926), .ZN(
        n5904) );
  OAI22_X1 U14286 ( .A1(n17132), .A2(n17443), .B1(n17129), .B2(n12925), .ZN(
        n5905) );
  OAI22_X1 U14287 ( .A1(n17132), .A2(n17445), .B1(n17129), .B2(n12924), .ZN(
        n5906) );
  OAI22_X1 U14288 ( .A1(n17132), .A2(n17447), .B1(n17129), .B2(n12923), .ZN(
        n5907) );
  OAI22_X1 U14289 ( .A1(n17132), .A2(n17449), .B1(n17129), .B2(n12922), .ZN(
        n5908) );
  OAI22_X1 U14290 ( .A1(n17132), .A2(n17451), .B1(n17129), .B2(n12921), .ZN(
        n5909) );
  OAI22_X1 U14291 ( .A1(n17133), .A2(n17453), .B1(n17129), .B2(n12920), .ZN(
        n5910) );
  OAI22_X1 U14292 ( .A1(n17133), .A2(n17455), .B1(n17129), .B2(n12919), .ZN(
        n5911) );
  OAI22_X1 U14293 ( .A1(n17133), .A2(n17457), .B1(n17130), .B2(n12918), .ZN(
        n5912) );
  OAI22_X1 U14294 ( .A1(n17133), .A2(n17459), .B1(n17130), .B2(n12917), .ZN(
        n5913) );
  OAI22_X1 U14295 ( .A1(n17133), .A2(n17461), .B1(n17130), .B2(n12916), .ZN(
        n5914) );
  OAI22_X1 U14296 ( .A1(n17134), .A2(n17463), .B1(n17130), .B2(n12915), .ZN(
        n5915) );
  OAI22_X1 U14297 ( .A1(n17134), .A2(n17465), .B1(n17130), .B2(n12914), .ZN(
        n5916) );
  OAI22_X1 U14298 ( .A1(n17134), .A2(n17467), .B1(n17130), .B2(n12913), .ZN(
        n5917) );
  OAI22_X1 U14299 ( .A1(n17134), .A2(n17469), .B1(n17130), .B2(n12912), .ZN(
        n5918) );
  OAI22_X1 U14300 ( .A1(n17134), .A2(n17471), .B1(n17130), .B2(n12911), .ZN(
        n5919) );
  OAI22_X1 U14301 ( .A1(n17135), .A2(n17473), .B1(n17130), .B2(n12910), .ZN(
        n5920) );
  OAI22_X1 U14302 ( .A1(n17135), .A2(n17475), .B1(n17130), .B2(n12909), .ZN(
        n5921) );
  OAI22_X1 U14303 ( .A1(n17135), .A2(n17477), .B1(n17130), .B2(n12908), .ZN(
        n5922) );
  OAI22_X1 U14304 ( .A1(n17135), .A2(n17479), .B1(n17130), .B2(n12907), .ZN(
        n5923) );
  OAI22_X1 U14305 ( .A1(n17148), .A2(n17433), .B1(n17146), .B2(n12866), .ZN(
        n5964) );
  OAI22_X1 U14306 ( .A1(n17148), .A2(n17435), .B1(n17146), .B2(n12865), .ZN(
        n5965) );
  OAI22_X1 U14307 ( .A1(n17148), .A2(n17437), .B1(n17146), .B2(n12864), .ZN(
        n5966) );
  OAI22_X1 U14308 ( .A1(n17148), .A2(n17439), .B1(n17146), .B2(n12863), .ZN(
        n5967) );
  OAI22_X1 U14309 ( .A1(n17148), .A2(n17441), .B1(n17146), .B2(n12862), .ZN(
        n5968) );
  OAI22_X1 U14310 ( .A1(n17149), .A2(n17443), .B1(n17146), .B2(n12861), .ZN(
        n5969) );
  OAI22_X1 U14311 ( .A1(n17149), .A2(n17445), .B1(n17146), .B2(n12860), .ZN(
        n5970) );
  OAI22_X1 U14312 ( .A1(n17149), .A2(n17447), .B1(n17146), .B2(n12859), .ZN(
        n5971) );
  OAI22_X1 U14313 ( .A1(n17149), .A2(n17449), .B1(n17146), .B2(n12858), .ZN(
        n5972) );
  OAI22_X1 U14314 ( .A1(n17149), .A2(n17451), .B1(n17146), .B2(n12857), .ZN(
        n5973) );
  OAI22_X1 U14315 ( .A1(n17150), .A2(n17453), .B1(n17146), .B2(n12856), .ZN(
        n5974) );
  OAI22_X1 U14316 ( .A1(n17150), .A2(n17455), .B1(n17146), .B2(n12855), .ZN(
        n5975) );
  OAI22_X1 U14317 ( .A1(n17150), .A2(n17457), .B1(n17147), .B2(n12854), .ZN(
        n5976) );
  OAI22_X1 U14318 ( .A1(n17150), .A2(n17459), .B1(n17147), .B2(n12853), .ZN(
        n5977) );
  OAI22_X1 U14319 ( .A1(n17150), .A2(n17461), .B1(n17147), .B2(n12852), .ZN(
        n5978) );
  OAI22_X1 U14320 ( .A1(n17151), .A2(n17463), .B1(n17147), .B2(n12851), .ZN(
        n5979) );
  OAI22_X1 U14321 ( .A1(n17151), .A2(n17465), .B1(n17147), .B2(n12850), .ZN(
        n5980) );
  OAI22_X1 U14322 ( .A1(n17151), .A2(n17467), .B1(n17147), .B2(n12849), .ZN(
        n5981) );
  OAI22_X1 U14323 ( .A1(n17151), .A2(n17469), .B1(n17147), .B2(n12848), .ZN(
        n5982) );
  OAI22_X1 U14324 ( .A1(n17151), .A2(n17471), .B1(n17147), .B2(n12847), .ZN(
        n5983) );
  OAI22_X1 U14325 ( .A1(n17152), .A2(n17473), .B1(n17147), .B2(n12846), .ZN(
        n5984) );
  OAI22_X1 U14326 ( .A1(n17152), .A2(n17475), .B1(n17147), .B2(n12845), .ZN(
        n5985) );
  OAI22_X1 U14327 ( .A1(n17152), .A2(n17477), .B1(n17147), .B2(n12844), .ZN(
        n5986) );
  OAI22_X1 U14328 ( .A1(n17152), .A2(n17479), .B1(n17147), .B2(n12843), .ZN(
        n5987) );
  OAI22_X1 U14329 ( .A1(n17268), .A2(n17433), .B1(n17266), .B2(n12581), .ZN(
        n6412) );
  OAI22_X1 U14330 ( .A1(n17268), .A2(n17435), .B1(n17266), .B2(n12580), .ZN(
        n6413) );
  OAI22_X1 U14331 ( .A1(n17268), .A2(n17437), .B1(n17266), .B2(n12579), .ZN(
        n6414) );
  OAI22_X1 U14332 ( .A1(n17268), .A2(n17439), .B1(n17266), .B2(n12578), .ZN(
        n6415) );
  OAI22_X1 U14333 ( .A1(n17268), .A2(n17441), .B1(n17266), .B2(n12577), .ZN(
        n6416) );
  OAI22_X1 U14334 ( .A1(n17269), .A2(n17443), .B1(n17266), .B2(n12576), .ZN(
        n6417) );
  OAI22_X1 U14335 ( .A1(n17269), .A2(n17445), .B1(n17266), .B2(n12575), .ZN(
        n6418) );
  OAI22_X1 U14336 ( .A1(n17269), .A2(n17447), .B1(n17266), .B2(n12574), .ZN(
        n6419) );
  OAI22_X1 U14337 ( .A1(n17269), .A2(n17449), .B1(n17266), .B2(n12573), .ZN(
        n6420) );
  OAI22_X1 U14338 ( .A1(n17269), .A2(n17451), .B1(n17266), .B2(n12572), .ZN(
        n6421) );
  OAI22_X1 U14339 ( .A1(n17270), .A2(n17453), .B1(n17266), .B2(n12571), .ZN(
        n6422) );
  OAI22_X1 U14340 ( .A1(n17270), .A2(n17455), .B1(n17266), .B2(n12570), .ZN(
        n6423) );
  OAI22_X1 U14341 ( .A1(n17270), .A2(n17457), .B1(n17267), .B2(n12569), .ZN(
        n6424) );
  OAI22_X1 U14342 ( .A1(n17270), .A2(n17459), .B1(n17267), .B2(n12568), .ZN(
        n6425) );
  OAI22_X1 U14343 ( .A1(n17270), .A2(n17461), .B1(n17267), .B2(n12567), .ZN(
        n6426) );
  OAI22_X1 U14344 ( .A1(n17271), .A2(n17463), .B1(n17267), .B2(n12566), .ZN(
        n6427) );
  OAI22_X1 U14345 ( .A1(n17271), .A2(n17465), .B1(n17267), .B2(n12565), .ZN(
        n6428) );
  OAI22_X1 U14346 ( .A1(n17271), .A2(n17467), .B1(n17267), .B2(n12564), .ZN(
        n6429) );
  OAI22_X1 U14347 ( .A1(n17271), .A2(n17469), .B1(n17267), .B2(n12563), .ZN(
        n6430) );
  OAI22_X1 U14348 ( .A1(n17271), .A2(n17471), .B1(n17267), .B2(n12562), .ZN(
        n6431) );
  OAI22_X1 U14349 ( .A1(n17272), .A2(n17473), .B1(n17267), .B2(n12561), .ZN(
        n6432) );
  OAI22_X1 U14350 ( .A1(n17272), .A2(n17475), .B1(n17267), .B2(n12560), .ZN(
        n6433) );
  OAI22_X1 U14351 ( .A1(n17272), .A2(n17477), .B1(n17267), .B2(n12559), .ZN(
        n6434) );
  OAI22_X1 U14352 ( .A1(n17272), .A2(n17479), .B1(n17267), .B2(n12558), .ZN(
        n6435) );
  OAI22_X1 U14353 ( .A1(n17285), .A2(n17433), .B1(n17283), .B2(n12517), .ZN(
        n6476) );
  OAI22_X1 U14354 ( .A1(n17285), .A2(n17435), .B1(n17283), .B2(n12516), .ZN(
        n6477) );
  OAI22_X1 U14355 ( .A1(n17285), .A2(n17437), .B1(n17283), .B2(n12515), .ZN(
        n6478) );
  OAI22_X1 U14356 ( .A1(n17285), .A2(n17439), .B1(n17283), .B2(n12514), .ZN(
        n6479) );
  OAI22_X1 U14357 ( .A1(n17285), .A2(n17441), .B1(n17283), .B2(n12513), .ZN(
        n6480) );
  OAI22_X1 U14358 ( .A1(n17286), .A2(n17443), .B1(n17283), .B2(n12512), .ZN(
        n6481) );
  OAI22_X1 U14359 ( .A1(n17286), .A2(n17445), .B1(n17283), .B2(n12511), .ZN(
        n6482) );
  OAI22_X1 U14360 ( .A1(n17286), .A2(n17447), .B1(n17283), .B2(n12510), .ZN(
        n6483) );
  OAI22_X1 U14361 ( .A1(n17286), .A2(n17449), .B1(n17283), .B2(n12509), .ZN(
        n6484) );
  OAI22_X1 U14362 ( .A1(n17286), .A2(n17451), .B1(n17283), .B2(n12508), .ZN(
        n6485) );
  OAI22_X1 U14363 ( .A1(n17287), .A2(n17453), .B1(n17283), .B2(n12507), .ZN(
        n6486) );
  OAI22_X1 U14364 ( .A1(n17287), .A2(n17455), .B1(n17283), .B2(n12506), .ZN(
        n6487) );
  OAI22_X1 U14365 ( .A1(n17287), .A2(n17457), .B1(n17284), .B2(n12505), .ZN(
        n6488) );
  OAI22_X1 U14366 ( .A1(n17287), .A2(n17459), .B1(n17284), .B2(n12504), .ZN(
        n6489) );
  OAI22_X1 U14367 ( .A1(n17287), .A2(n17461), .B1(n17284), .B2(n12503), .ZN(
        n6490) );
  OAI22_X1 U14368 ( .A1(n17288), .A2(n17463), .B1(n17284), .B2(n12502), .ZN(
        n6491) );
  OAI22_X1 U14369 ( .A1(n17288), .A2(n17465), .B1(n17284), .B2(n12501), .ZN(
        n6492) );
  OAI22_X1 U14370 ( .A1(n17288), .A2(n17467), .B1(n17284), .B2(n12500), .ZN(
        n6493) );
  OAI22_X1 U14371 ( .A1(n17288), .A2(n17469), .B1(n17284), .B2(n12499), .ZN(
        n6494) );
  OAI22_X1 U14372 ( .A1(n17288), .A2(n17471), .B1(n17284), .B2(n12498), .ZN(
        n6495) );
  OAI22_X1 U14373 ( .A1(n17289), .A2(n17473), .B1(n17284), .B2(n12497), .ZN(
        n6496) );
  OAI22_X1 U14374 ( .A1(n17289), .A2(n17475), .B1(n17284), .B2(n12496), .ZN(
        n6497) );
  OAI22_X1 U14375 ( .A1(n17289), .A2(n17477), .B1(n17284), .B2(n12495), .ZN(
        n6498) );
  OAI22_X1 U14376 ( .A1(n17289), .A2(n17479), .B1(n17284), .B2(n12494), .ZN(
        n6499) );
  OAI221_X1 U14377 ( .B1(n7864), .B2(n16631), .C1(n8055), .C2(n16625), .A(
        n16075), .ZN(n16059) );
  AOI22_X1 U14378 ( .A1(n16619), .A2(n13186), .B1(n16613), .B2(n8120), .ZN(
        n16075) );
  OAI221_X1 U14379 ( .B1(n16413), .B2(n16577), .C1(n16414), .C2(n16571), .A(
        n16081), .ZN(n16080) );
  AOI22_X1 U14380 ( .A1(n16565), .A2(n12389), .B1(n16560), .B2(OUT2[0]), .ZN(
        n16081) );
  OAI221_X1 U14381 ( .B1(n7862), .B2(n16631), .C1(n8052), .C2(n16625), .A(
        n16046), .ZN(n16041) );
  AOI22_X1 U14382 ( .A1(n16619), .A2(n13185), .B1(n16613), .B2(n8119), .ZN(
        n16046) );
  OAI221_X1 U14383 ( .B1(n16408), .B2(n16577), .C1(n16409), .C2(n16571), .A(
        n16052), .ZN(n16051) );
  AOI22_X1 U14384 ( .A1(n16565), .A2(n12388), .B1(n16560), .B2(OUT2[1]), .ZN(
        n16052) );
  OAI221_X1 U14385 ( .B1(n7860), .B2(n16631), .C1(n8049), .C2(n16625), .A(
        n16028), .ZN(n16023) );
  AOI22_X1 U14386 ( .A1(n16619), .A2(n13184), .B1(n16613), .B2(n8118), .ZN(
        n16028) );
  OAI221_X1 U14387 ( .B1(n16403), .B2(n16577), .C1(n16404), .C2(n16571), .A(
        n16034), .ZN(n16033) );
  AOI22_X1 U14388 ( .A1(n16565), .A2(n12387), .B1(n16560), .B2(OUT2[2]), .ZN(
        n16034) );
  OAI221_X1 U14389 ( .B1(n7858), .B2(n16631), .C1(n8046), .C2(n16625), .A(
        n16010), .ZN(n16005) );
  AOI22_X1 U14390 ( .A1(n16619), .A2(n13183), .B1(n16613), .B2(n8117), .ZN(
        n16010) );
  OAI221_X1 U14391 ( .B1(n16398), .B2(n16577), .C1(n16399), .C2(n16571), .A(
        n16016), .ZN(n16015) );
  AOI22_X1 U14392 ( .A1(n16565), .A2(n12386), .B1(n16560), .B2(OUT2[3]), .ZN(
        n16016) );
  OAI221_X1 U14393 ( .B1(n7856), .B2(n16631), .C1(n8043), .C2(n16625), .A(
        n15992), .ZN(n15987) );
  AOI22_X1 U14394 ( .A1(n16619), .A2(n13182), .B1(n16613), .B2(n8116), .ZN(
        n15992) );
  OAI221_X1 U14395 ( .B1(n16393), .B2(n16577), .C1(n16394), .C2(n16571), .A(
        n15998), .ZN(n15997) );
  AOI22_X1 U14396 ( .A1(n16565), .A2(n12385), .B1(n16560), .B2(OUT2[4]), .ZN(
        n15998) );
  OAI221_X1 U14397 ( .B1(n7854), .B2(n16631), .C1(n8040), .C2(n16625), .A(
        n15974), .ZN(n15969) );
  AOI22_X1 U14398 ( .A1(n16619), .A2(n13181), .B1(n16613), .B2(n8115), .ZN(
        n15974) );
  OAI221_X1 U14399 ( .B1(n16388), .B2(n16577), .C1(n16389), .C2(n16571), .A(
        n15980), .ZN(n15979) );
  AOI22_X1 U14400 ( .A1(n16565), .A2(n12384), .B1(n16560), .B2(OUT2[5]), .ZN(
        n15980) );
  OAI221_X1 U14401 ( .B1(n7852), .B2(n16631), .C1(n8037), .C2(n16625), .A(
        n15956), .ZN(n15951) );
  AOI22_X1 U14402 ( .A1(n16619), .A2(n13180), .B1(n16613), .B2(n8114), .ZN(
        n15956) );
  OAI221_X1 U14403 ( .B1(n16383), .B2(n16577), .C1(n16384), .C2(n16571), .A(
        n15962), .ZN(n15961) );
  AOI22_X1 U14404 ( .A1(n16565), .A2(n12383), .B1(n16560), .B2(OUT2[6]), .ZN(
        n15962) );
  OAI221_X1 U14405 ( .B1(n7850), .B2(n16631), .C1(n8034), .C2(n16625), .A(
        n15938), .ZN(n15933) );
  AOI22_X1 U14406 ( .A1(n16619), .A2(n13179), .B1(n16613), .B2(n8113), .ZN(
        n15938) );
  OAI221_X1 U14407 ( .B1(n16378), .B2(n16577), .C1(n16379), .C2(n16571), .A(
        n15944), .ZN(n15943) );
  AOI22_X1 U14408 ( .A1(n16565), .A2(n12382), .B1(n16560), .B2(OUT2[7]), .ZN(
        n15944) );
  OAI221_X1 U14409 ( .B1(n7848), .B2(n16631), .C1(n8031), .C2(n16625), .A(
        n15920), .ZN(n15915) );
  AOI22_X1 U14410 ( .A1(n16619), .A2(n13178), .B1(n16613), .B2(n8112), .ZN(
        n15920) );
  OAI221_X1 U14411 ( .B1(n16373), .B2(n16577), .C1(n16374), .C2(n16571), .A(
        n15926), .ZN(n15925) );
  AOI22_X1 U14412 ( .A1(n16565), .A2(n12381), .B1(n16560), .B2(OUT2[8]), .ZN(
        n15926) );
  OAI221_X1 U14413 ( .B1(n7846), .B2(n16631), .C1(n8028), .C2(n16625), .A(
        n15902), .ZN(n15897) );
  AOI22_X1 U14414 ( .A1(n16619), .A2(n13177), .B1(n16613), .B2(n8111), .ZN(
        n15902) );
  OAI221_X1 U14415 ( .B1(n16368), .B2(n16577), .C1(n16369), .C2(n16571), .A(
        n15908), .ZN(n15907) );
  AOI22_X1 U14416 ( .A1(n16565), .A2(n12380), .B1(n16560), .B2(OUT2[9]), .ZN(
        n15908) );
  OAI221_X1 U14417 ( .B1(n7844), .B2(n16631), .C1(n8025), .C2(n16625), .A(
        n15884), .ZN(n15879) );
  AOI22_X1 U14418 ( .A1(n16619), .A2(n13176), .B1(n16613), .B2(n8110), .ZN(
        n15884) );
  OAI221_X1 U14419 ( .B1(n16363), .B2(n16577), .C1(n16364), .C2(n16571), .A(
        n15890), .ZN(n15889) );
  AOI22_X1 U14420 ( .A1(n16565), .A2(n12379), .B1(n16560), .B2(OUT2[10]), .ZN(
        n15890) );
  OAI221_X1 U14421 ( .B1(n7842), .B2(n16631), .C1(n8022), .C2(n16625), .A(
        n15866), .ZN(n15861) );
  AOI22_X1 U14422 ( .A1(n16619), .A2(n13175), .B1(n16613), .B2(n8109), .ZN(
        n15866) );
  OAI221_X1 U14423 ( .B1(n16358), .B2(n16577), .C1(n16359), .C2(n16571), .A(
        n15872), .ZN(n15871) );
  AOI22_X1 U14424 ( .A1(n16565), .A2(n12378), .B1(n16561), .B2(OUT2[11]), .ZN(
        n15872) );
  OAI221_X1 U14425 ( .B1(n7840), .B2(n16632), .C1(n8019), .C2(n16626), .A(
        n15848), .ZN(n15843) );
  AOI22_X1 U14426 ( .A1(n16620), .A2(n13174), .B1(n16614), .B2(n8108), .ZN(
        n15848) );
  OAI221_X1 U14427 ( .B1(n16353), .B2(n16578), .C1(n16354), .C2(n16572), .A(
        n15854), .ZN(n15853) );
  AOI22_X1 U14428 ( .A1(n16566), .A2(n12377), .B1(n16561), .B2(OUT2[12]), .ZN(
        n15854) );
  OAI221_X1 U14429 ( .B1(n7838), .B2(n16632), .C1(n8016), .C2(n16626), .A(
        n15830), .ZN(n15825) );
  AOI22_X1 U14430 ( .A1(n16620), .A2(n13173), .B1(n16614), .B2(n8107), .ZN(
        n15830) );
  OAI221_X1 U14431 ( .B1(n16348), .B2(n16578), .C1(n16349), .C2(n16572), .A(
        n15836), .ZN(n15835) );
  AOI22_X1 U14432 ( .A1(n16566), .A2(n12376), .B1(n16561), .B2(OUT2[13]), .ZN(
        n15836) );
  OAI221_X1 U14433 ( .B1(n7836), .B2(n16632), .C1(n8013), .C2(n16626), .A(
        n15812), .ZN(n15807) );
  AOI22_X1 U14434 ( .A1(n16620), .A2(n13172), .B1(n16614), .B2(n8106), .ZN(
        n15812) );
  OAI221_X1 U14435 ( .B1(n16343), .B2(n16578), .C1(n16344), .C2(n16572), .A(
        n15818), .ZN(n15817) );
  AOI22_X1 U14436 ( .A1(n16566), .A2(n12375), .B1(n16561), .B2(OUT2[14]), .ZN(
        n15818) );
  OAI221_X1 U14437 ( .B1(n7834), .B2(n16632), .C1(n8010), .C2(n16626), .A(
        n15794), .ZN(n15789) );
  AOI22_X1 U14438 ( .A1(n16620), .A2(n13171), .B1(n16614), .B2(n8105), .ZN(
        n15794) );
  OAI221_X1 U14439 ( .B1(n16338), .B2(n16578), .C1(n16339), .C2(n16572), .A(
        n15800), .ZN(n15799) );
  AOI22_X1 U14440 ( .A1(n16566), .A2(n12374), .B1(n16561), .B2(OUT2[15]), .ZN(
        n15800) );
  OAI221_X1 U14441 ( .B1(n7832), .B2(n16632), .C1(n8007), .C2(n16626), .A(
        n15776), .ZN(n15771) );
  AOI22_X1 U14442 ( .A1(n16620), .A2(n13170), .B1(n16614), .B2(n8104), .ZN(
        n15776) );
  OAI221_X1 U14443 ( .B1(n16333), .B2(n16578), .C1(n16334), .C2(n16572), .A(
        n15782), .ZN(n15781) );
  AOI22_X1 U14444 ( .A1(n16566), .A2(n12373), .B1(n16561), .B2(OUT2[16]), .ZN(
        n15782) );
  OAI221_X1 U14445 ( .B1(n7830), .B2(n16632), .C1(n8004), .C2(n16626), .A(
        n15758), .ZN(n15753) );
  AOI22_X1 U14446 ( .A1(n16620), .A2(n13169), .B1(n16614), .B2(n8103), .ZN(
        n15758) );
  OAI221_X1 U14447 ( .B1(n16328), .B2(n16578), .C1(n16329), .C2(n16572), .A(
        n15764), .ZN(n15763) );
  AOI22_X1 U14448 ( .A1(n16566), .A2(n12372), .B1(n16561), .B2(OUT2[17]), .ZN(
        n15764) );
  OAI221_X1 U14449 ( .B1(n7828), .B2(n16632), .C1(n8001), .C2(n16626), .A(
        n15740), .ZN(n15735) );
  AOI22_X1 U14450 ( .A1(n16620), .A2(n13168), .B1(n16614), .B2(n8102), .ZN(
        n15740) );
  OAI221_X1 U14451 ( .B1(n16323), .B2(n16578), .C1(n16324), .C2(n16572), .A(
        n15746), .ZN(n15745) );
  AOI22_X1 U14452 ( .A1(n16566), .A2(n12371), .B1(n16561), .B2(OUT2[18]), .ZN(
        n15746) );
  OAI221_X1 U14453 ( .B1(n7826), .B2(n16632), .C1(n7998), .C2(n16626), .A(
        n15722), .ZN(n15717) );
  AOI22_X1 U14454 ( .A1(n16620), .A2(n13167), .B1(n16614), .B2(n8101), .ZN(
        n15722) );
  OAI221_X1 U14455 ( .B1(n16318), .B2(n16578), .C1(n16319), .C2(n16572), .A(
        n15728), .ZN(n15727) );
  AOI22_X1 U14456 ( .A1(n16566), .A2(n12370), .B1(n16561), .B2(OUT2[19]), .ZN(
        n15728) );
  OAI221_X1 U14457 ( .B1(n7824), .B2(n16632), .C1(n7995), .C2(n16626), .A(
        n15704), .ZN(n15699) );
  AOI22_X1 U14458 ( .A1(n16620), .A2(n13166), .B1(n16614), .B2(n8100), .ZN(
        n15704) );
  OAI221_X1 U14459 ( .B1(n16313), .B2(n16578), .C1(n16314), .C2(n16572), .A(
        n15710), .ZN(n15709) );
  AOI22_X1 U14460 ( .A1(n16566), .A2(n12369), .B1(n16561), .B2(OUT2[20]), .ZN(
        n15710) );
  OAI221_X1 U14461 ( .B1(n7822), .B2(n16632), .C1(n7992), .C2(n16626), .A(
        n15686), .ZN(n15681) );
  AOI22_X1 U14462 ( .A1(n16620), .A2(n13165), .B1(n16614), .B2(n8099), .ZN(
        n15686) );
  OAI221_X1 U14463 ( .B1(n16308), .B2(n16578), .C1(n16309), .C2(n16572), .A(
        n15692), .ZN(n15691) );
  AOI22_X1 U14464 ( .A1(n16566), .A2(n12368), .B1(n16561), .B2(OUT2[21]), .ZN(
        n15692) );
  OAI221_X1 U14465 ( .B1(n7820), .B2(n16632), .C1(n7989), .C2(n16626), .A(
        n15668), .ZN(n15663) );
  AOI22_X1 U14466 ( .A1(n16620), .A2(n13164), .B1(n16614), .B2(n8098), .ZN(
        n15668) );
  OAI221_X1 U14467 ( .B1(n16303), .B2(n16578), .C1(n16304), .C2(n16572), .A(
        n15674), .ZN(n15673) );
  AOI22_X1 U14468 ( .A1(n16566), .A2(n12367), .B1(n16561), .B2(OUT2[22]), .ZN(
        n15674) );
  OAI221_X1 U14469 ( .B1(n7818), .B2(n16632), .C1(n7986), .C2(n16626), .A(
        n15650), .ZN(n15645) );
  AOI22_X1 U14470 ( .A1(n16620), .A2(n13163), .B1(n16614), .B2(n8097), .ZN(
        n15650) );
  OAI221_X1 U14471 ( .B1(n16298), .B2(n16578), .C1(n16299), .C2(n16572), .A(
        n15656), .ZN(n15655) );
  AOI22_X1 U14472 ( .A1(n16566), .A2(n12366), .B1(n16561), .B2(OUT2[23]), .ZN(
        n15656) );
  OAI221_X1 U14473 ( .B1(n7816), .B2(n16633), .C1(n7983), .C2(n16627), .A(
        n15632), .ZN(n15627) );
  AOI22_X1 U14474 ( .A1(n16621), .A2(n13162), .B1(n16615), .B2(n8096), .ZN(
        n15632) );
  OAI221_X1 U14475 ( .B1(n16293), .B2(n16579), .C1(n16294), .C2(n16573), .A(
        n15638), .ZN(n15637) );
  AOI22_X1 U14476 ( .A1(n16567), .A2(n12365), .B1(n16562), .B2(OUT2[24]), .ZN(
        n15638) );
  OAI221_X1 U14477 ( .B1(n7814), .B2(n16633), .C1(n7980), .C2(n16627), .A(
        n15614), .ZN(n15609) );
  AOI22_X1 U14478 ( .A1(n16621), .A2(n13161), .B1(n16615), .B2(n8095), .ZN(
        n15614) );
  OAI221_X1 U14479 ( .B1(n16288), .B2(n16579), .C1(n16289), .C2(n16573), .A(
        n15620), .ZN(n15619) );
  AOI22_X1 U14480 ( .A1(n16567), .A2(n12364), .B1(n16562), .B2(OUT2[25]), .ZN(
        n15620) );
  OAI221_X1 U14481 ( .B1(n7812), .B2(n16633), .C1(n7977), .C2(n16627), .A(
        n15596), .ZN(n15591) );
  AOI22_X1 U14482 ( .A1(n16621), .A2(n13160), .B1(n16615), .B2(n8094), .ZN(
        n15596) );
  OAI221_X1 U14483 ( .B1(n16283), .B2(n16579), .C1(n16284), .C2(n16573), .A(
        n15602), .ZN(n15601) );
  AOI22_X1 U14484 ( .A1(n16567), .A2(n12363), .B1(n16562), .B2(OUT2[26]), .ZN(
        n15602) );
  OAI221_X1 U14485 ( .B1(n7810), .B2(n16633), .C1(n7974), .C2(n16627), .A(
        n15578), .ZN(n15573) );
  AOI22_X1 U14486 ( .A1(n16621), .A2(n13159), .B1(n16615), .B2(n8093), .ZN(
        n15578) );
  OAI221_X1 U14487 ( .B1(n16278), .B2(n16579), .C1(n16279), .C2(n16573), .A(
        n15584), .ZN(n15583) );
  AOI22_X1 U14488 ( .A1(n16567), .A2(n12362), .B1(n16562), .B2(OUT2[27]), .ZN(
        n15584) );
  OAI221_X1 U14489 ( .B1(n7808), .B2(n16633), .C1(n7971), .C2(n16627), .A(
        n15560), .ZN(n15555) );
  AOI22_X1 U14490 ( .A1(n16621), .A2(n13158), .B1(n16615), .B2(n8092), .ZN(
        n15560) );
  OAI221_X1 U14491 ( .B1(n16273), .B2(n16579), .C1(n16274), .C2(n16573), .A(
        n15566), .ZN(n15565) );
  AOI22_X1 U14492 ( .A1(n16567), .A2(n12361), .B1(n16562), .B2(OUT2[28]), .ZN(
        n15566) );
  OAI221_X1 U14493 ( .B1(n7806), .B2(n16633), .C1(n7968), .C2(n16627), .A(
        n15542), .ZN(n15537) );
  AOI22_X1 U14494 ( .A1(n16621), .A2(n13157), .B1(n16615), .B2(n8091), .ZN(
        n15542) );
  OAI221_X1 U14495 ( .B1(n16268), .B2(n16579), .C1(n16269), .C2(n16573), .A(
        n15548), .ZN(n15547) );
  AOI22_X1 U14496 ( .A1(n16567), .A2(n12360), .B1(n16562), .B2(OUT2[29]), .ZN(
        n15548) );
  OAI221_X1 U14497 ( .B1(n7804), .B2(n16633), .C1(n7965), .C2(n16627), .A(
        n15524), .ZN(n15519) );
  AOI22_X1 U14498 ( .A1(n16621), .A2(n13156), .B1(n16615), .B2(n8090), .ZN(
        n15524) );
  OAI221_X1 U14499 ( .B1(n16263), .B2(n16579), .C1(n16264), .C2(n16573), .A(
        n15530), .ZN(n15529) );
  AOI22_X1 U14500 ( .A1(n16567), .A2(n12359), .B1(n16562), .B2(OUT2[30]), .ZN(
        n15530) );
  OAI221_X1 U14501 ( .B1(n7802), .B2(n16633), .C1(n7962), .C2(n16627), .A(
        n15506), .ZN(n15501) );
  AOI22_X1 U14502 ( .A1(n16621), .A2(n13155), .B1(n16615), .B2(n8089), .ZN(
        n15506) );
  OAI221_X1 U14503 ( .B1(n16258), .B2(n16579), .C1(n16259), .C2(n16573), .A(
        n15512), .ZN(n15511) );
  AOI22_X1 U14504 ( .A1(n16567), .A2(n12358), .B1(n16562), .B2(OUT2[31]), .ZN(
        n15512) );
  OAI221_X1 U14505 ( .B1(n7800), .B2(n16633), .C1(n7959), .C2(n16627), .A(
        n15488), .ZN(n15483) );
  AOI22_X1 U14506 ( .A1(n16621), .A2(n13154), .B1(n16615), .B2(n8088), .ZN(
        n15488) );
  OAI221_X1 U14507 ( .B1(n16253), .B2(n16579), .C1(n16254), .C2(n16573), .A(
        n15494), .ZN(n15493) );
  AOI22_X1 U14508 ( .A1(n16567), .A2(n12357), .B1(n16562), .B2(OUT2[32]), .ZN(
        n15494) );
  OAI221_X1 U14509 ( .B1(n7798), .B2(n16633), .C1(n7956), .C2(n16627), .A(
        n15470), .ZN(n15465) );
  AOI22_X1 U14510 ( .A1(n16621), .A2(n13153), .B1(n16615), .B2(n8087), .ZN(
        n15470) );
  OAI221_X1 U14511 ( .B1(n16248), .B2(n16579), .C1(n16249), .C2(n16573), .A(
        n15476), .ZN(n15475) );
  AOI22_X1 U14512 ( .A1(n16567), .A2(n12356), .B1(n16562), .B2(OUT2[33]), .ZN(
        n15476) );
  OAI221_X1 U14513 ( .B1(n7796), .B2(n16633), .C1(n7953), .C2(n16627), .A(
        n15452), .ZN(n15447) );
  AOI22_X1 U14514 ( .A1(n16621), .A2(n13152), .B1(n16615), .B2(n8086), .ZN(
        n15452) );
  OAI221_X1 U14515 ( .B1(n16243), .B2(n16579), .C1(n16244), .C2(n16573), .A(
        n15458), .ZN(n15457) );
  AOI22_X1 U14516 ( .A1(n16567), .A2(n12355), .B1(n16562), .B2(OUT2[34]), .ZN(
        n15458) );
  OAI221_X1 U14517 ( .B1(n7794), .B2(n16633), .C1(n7950), .C2(n16627), .A(
        n15434), .ZN(n15429) );
  AOI22_X1 U14518 ( .A1(n16621), .A2(n13151), .B1(n16615), .B2(n8085), .ZN(
        n15434) );
  OAI221_X1 U14519 ( .B1(n16238), .B2(n16579), .C1(n16239), .C2(n16573), .A(
        n15440), .ZN(n15439) );
  AOI22_X1 U14520 ( .A1(n16567), .A2(n12354), .B1(n16562), .B2(OUT2[35]), .ZN(
        n15440) );
  OAI221_X1 U14521 ( .B1(n7792), .B2(n16634), .C1(n7947), .C2(n16628), .A(
        n15416), .ZN(n15411) );
  AOI22_X1 U14522 ( .A1(n16622), .A2(n13150), .B1(n16616), .B2(n8084), .ZN(
        n15416) );
  OAI221_X1 U14523 ( .B1(n16233), .B2(n16580), .C1(n16234), .C2(n16574), .A(
        n15422), .ZN(n15421) );
  AOI22_X1 U14524 ( .A1(n16568), .A2(n12353), .B1(n16562), .B2(OUT2[36]), .ZN(
        n15422) );
  OAI221_X1 U14525 ( .B1(n7790), .B2(n16634), .C1(n7944), .C2(n16628), .A(
        n15398), .ZN(n15393) );
  AOI22_X1 U14526 ( .A1(n16622), .A2(n13149), .B1(n16616), .B2(n8083), .ZN(
        n15398) );
  OAI221_X1 U14527 ( .B1(n16228), .B2(n16580), .C1(n16229), .C2(n16574), .A(
        n15404), .ZN(n15403) );
  AOI22_X1 U14528 ( .A1(n16568), .A2(n12352), .B1(n16563), .B2(OUT2[37]), .ZN(
        n15404) );
  OAI221_X1 U14529 ( .B1(n7788), .B2(n16634), .C1(n7941), .C2(n16628), .A(
        n15380), .ZN(n15375) );
  AOI22_X1 U14530 ( .A1(n16622), .A2(n13148), .B1(n16616), .B2(n8082), .ZN(
        n15380) );
  OAI221_X1 U14531 ( .B1(n16223), .B2(n16580), .C1(n16224), .C2(n16574), .A(
        n15386), .ZN(n15385) );
  AOI22_X1 U14532 ( .A1(n16568), .A2(n12351), .B1(n16563), .B2(OUT2[38]), .ZN(
        n15386) );
  OAI221_X1 U14533 ( .B1(n7786), .B2(n16634), .C1(n7938), .C2(n16628), .A(
        n15362), .ZN(n15357) );
  AOI22_X1 U14534 ( .A1(n16622), .A2(n13147), .B1(n16616), .B2(n8081), .ZN(
        n15362) );
  OAI221_X1 U14535 ( .B1(n16218), .B2(n16580), .C1(n16219), .C2(n16574), .A(
        n15368), .ZN(n15367) );
  AOI22_X1 U14536 ( .A1(n16568), .A2(n12350), .B1(n16563), .B2(OUT2[39]), .ZN(
        n15368) );
  OAI221_X1 U14537 ( .B1(n7784), .B2(n16634), .C1(n7935), .C2(n16628), .A(
        n15344), .ZN(n15339) );
  AOI22_X1 U14538 ( .A1(n16622), .A2(n13146), .B1(n16616), .B2(n8080), .ZN(
        n15344) );
  OAI221_X1 U14539 ( .B1(n16213), .B2(n16580), .C1(n16214), .C2(n16574), .A(
        n15350), .ZN(n15349) );
  AOI22_X1 U14540 ( .A1(n16568), .A2(n12349), .B1(n16563), .B2(OUT2[40]), .ZN(
        n15350) );
  OAI221_X1 U14541 ( .B1(n7782), .B2(n16634), .C1(n7932), .C2(n16628), .A(
        n15326), .ZN(n15321) );
  AOI22_X1 U14542 ( .A1(n16622), .A2(n13145), .B1(n16616), .B2(n8079), .ZN(
        n15326) );
  OAI221_X1 U14543 ( .B1(n16208), .B2(n16580), .C1(n16209), .C2(n16574), .A(
        n15332), .ZN(n15331) );
  AOI22_X1 U14544 ( .A1(n16568), .A2(n12348), .B1(n16563), .B2(OUT2[41]), .ZN(
        n15332) );
  OAI221_X1 U14545 ( .B1(n7780), .B2(n16634), .C1(n7929), .C2(n16628), .A(
        n15308), .ZN(n15303) );
  AOI22_X1 U14546 ( .A1(n16622), .A2(n13144), .B1(n16616), .B2(n8078), .ZN(
        n15308) );
  OAI221_X1 U14547 ( .B1(n16203), .B2(n16580), .C1(n16204), .C2(n16574), .A(
        n15314), .ZN(n15313) );
  AOI22_X1 U14548 ( .A1(n16568), .A2(n12347), .B1(n16563), .B2(OUT2[42]), .ZN(
        n15314) );
  OAI221_X1 U14549 ( .B1(n7778), .B2(n16634), .C1(n7926), .C2(n16628), .A(
        n15290), .ZN(n15285) );
  AOI22_X1 U14550 ( .A1(n16622), .A2(n13143), .B1(n16616), .B2(n8077), .ZN(
        n15290) );
  OAI221_X1 U14551 ( .B1(n16198), .B2(n16580), .C1(n16199), .C2(n16574), .A(
        n15296), .ZN(n15295) );
  AOI22_X1 U14552 ( .A1(n16568), .A2(n12346), .B1(n16563), .B2(OUT2[43]), .ZN(
        n15296) );
  OAI221_X1 U14553 ( .B1(n7776), .B2(n16634), .C1(n7923), .C2(n16628), .A(
        n15272), .ZN(n15267) );
  AOI22_X1 U14554 ( .A1(n16622), .A2(n13142), .B1(n16616), .B2(n8076), .ZN(
        n15272) );
  OAI221_X1 U14555 ( .B1(n16193), .B2(n16580), .C1(n16194), .C2(n16574), .A(
        n15278), .ZN(n15277) );
  AOI22_X1 U14556 ( .A1(n16568), .A2(n12345), .B1(n16563), .B2(OUT2[44]), .ZN(
        n15278) );
  OAI221_X1 U14557 ( .B1(n7774), .B2(n16634), .C1(n7920), .C2(n16628), .A(
        n15254), .ZN(n15249) );
  AOI22_X1 U14558 ( .A1(n16622), .A2(n13141), .B1(n16616), .B2(n8075), .ZN(
        n15254) );
  OAI221_X1 U14559 ( .B1(n16188), .B2(n16580), .C1(n16189), .C2(n16574), .A(
        n15260), .ZN(n15259) );
  AOI22_X1 U14560 ( .A1(n16568), .A2(n12344), .B1(n16563), .B2(OUT2[45]), .ZN(
        n15260) );
  OAI221_X1 U14561 ( .B1(n7772), .B2(n16634), .C1(n7917), .C2(n16628), .A(
        n15236), .ZN(n15231) );
  AOI22_X1 U14562 ( .A1(n16622), .A2(n13140), .B1(n16616), .B2(n8074), .ZN(
        n15236) );
  OAI221_X1 U14563 ( .B1(n16183), .B2(n16580), .C1(n16184), .C2(n16574), .A(
        n15242), .ZN(n15241) );
  AOI22_X1 U14564 ( .A1(n16568), .A2(n12343), .B1(n16563), .B2(OUT2[46]), .ZN(
        n15242) );
  OAI221_X1 U14565 ( .B1(n7770), .B2(n16634), .C1(n7914), .C2(n16628), .A(
        n15218), .ZN(n15213) );
  AOI22_X1 U14566 ( .A1(n16622), .A2(n13139), .B1(n16616), .B2(n8073), .ZN(
        n15218) );
  OAI221_X1 U14567 ( .B1(n16178), .B2(n16580), .C1(n16179), .C2(n16574), .A(
        n15224), .ZN(n15223) );
  AOI22_X1 U14568 ( .A1(n16568), .A2(n12342), .B1(n16563), .B2(OUT2[47]), .ZN(
        n15224) );
  OAI221_X1 U14569 ( .B1(n7768), .B2(n16635), .C1(n7911), .C2(n16629), .A(
        n15200), .ZN(n15195) );
  AOI22_X1 U14570 ( .A1(n16623), .A2(n13138), .B1(n16617), .B2(n8072), .ZN(
        n15200) );
  OAI221_X1 U14571 ( .B1(n16173), .B2(n16581), .C1(n16174), .C2(n16575), .A(
        n15206), .ZN(n15205) );
  AOI22_X1 U14572 ( .A1(n16569), .A2(n12341), .B1(n16563), .B2(OUT2[48]), .ZN(
        n15206) );
  OAI221_X1 U14573 ( .B1(n7766), .B2(n16635), .C1(n7908), .C2(n16629), .A(
        n15182), .ZN(n15177) );
  AOI22_X1 U14574 ( .A1(n16623), .A2(n13137), .B1(n16617), .B2(n8071), .ZN(
        n15182) );
  OAI221_X1 U14575 ( .B1(n16168), .B2(n16581), .C1(n16169), .C2(n16575), .A(
        n15188), .ZN(n15187) );
  AOI22_X1 U14576 ( .A1(n16569), .A2(n12340), .B1(n16563), .B2(OUT2[49]), .ZN(
        n15188) );
  OAI221_X1 U14577 ( .B1(n7764), .B2(n16635), .C1(n7905), .C2(n16629), .A(
        n15164), .ZN(n15159) );
  AOI22_X1 U14578 ( .A1(n16623), .A2(n13136), .B1(n16617), .B2(n8070), .ZN(
        n15164) );
  OAI221_X1 U14579 ( .B1(n16163), .B2(n16581), .C1(n16164), .C2(n16575), .A(
        n15170), .ZN(n15169) );
  AOI22_X1 U14580 ( .A1(n16569), .A2(n12339), .B1(n16564), .B2(OUT2[50]), .ZN(
        n15170) );
  OAI221_X1 U14581 ( .B1(n7762), .B2(n16635), .C1(n7902), .C2(n16629), .A(
        n15146), .ZN(n15141) );
  AOI22_X1 U14582 ( .A1(n16623), .A2(n13135), .B1(n16617), .B2(n8069), .ZN(
        n15146) );
  OAI221_X1 U14583 ( .B1(n16158), .B2(n16581), .C1(n16159), .C2(n16575), .A(
        n15152), .ZN(n15151) );
  AOI22_X1 U14584 ( .A1(n16569), .A2(n12338), .B1(n16564), .B2(OUT2[51]), .ZN(
        n15152) );
  OAI221_X1 U14585 ( .B1(n7760), .B2(n16635), .C1(n7899), .C2(n16629), .A(
        n15128), .ZN(n15123) );
  AOI22_X1 U14586 ( .A1(n16623), .A2(n13134), .B1(n16617), .B2(n8068), .ZN(
        n15128) );
  OAI221_X1 U14587 ( .B1(n16153), .B2(n16581), .C1(n16154), .C2(n16575), .A(
        n15134), .ZN(n15133) );
  AOI22_X1 U14588 ( .A1(n16569), .A2(n12337), .B1(n16564), .B2(OUT2[52]), .ZN(
        n15134) );
  OAI221_X1 U14589 ( .B1(n7758), .B2(n16635), .C1(n7896), .C2(n16629), .A(
        n15110), .ZN(n15105) );
  AOI22_X1 U14590 ( .A1(n16623), .A2(n13133), .B1(n16617), .B2(n8067), .ZN(
        n15110) );
  OAI221_X1 U14591 ( .B1(n16148), .B2(n16581), .C1(n16149), .C2(n16575), .A(
        n15116), .ZN(n15115) );
  AOI22_X1 U14592 ( .A1(n16569), .A2(n12336), .B1(n16564), .B2(OUT2[53]), .ZN(
        n15116) );
  OAI221_X1 U14593 ( .B1(n7756), .B2(n16635), .C1(n7893), .C2(n16629), .A(
        n15092), .ZN(n15087) );
  AOI22_X1 U14594 ( .A1(n16623), .A2(n13132), .B1(n16617), .B2(n8066), .ZN(
        n15092) );
  OAI221_X1 U14595 ( .B1(n16143), .B2(n16581), .C1(n16144), .C2(n16575), .A(
        n15098), .ZN(n15097) );
  AOI22_X1 U14596 ( .A1(n16569), .A2(n12335), .B1(n16564), .B2(OUT2[54]), .ZN(
        n15098) );
  OAI221_X1 U14597 ( .B1(n7754), .B2(n16635), .C1(n7890), .C2(n16629), .A(
        n15074), .ZN(n15069) );
  AOI22_X1 U14598 ( .A1(n16623), .A2(n13131), .B1(n16617), .B2(n8065), .ZN(
        n15074) );
  OAI221_X1 U14599 ( .B1(n16138), .B2(n16581), .C1(n16139), .C2(n16575), .A(
        n15080), .ZN(n15079) );
  AOI22_X1 U14600 ( .A1(n16569), .A2(n12334), .B1(n16564), .B2(OUT2[55]), .ZN(
        n15080) );
  OAI221_X1 U14601 ( .B1(n7752), .B2(n16635), .C1(n7887), .C2(n16629), .A(
        n15056), .ZN(n15051) );
  AOI22_X1 U14602 ( .A1(n16623), .A2(n13130), .B1(n16617), .B2(n8064), .ZN(
        n15056) );
  OAI221_X1 U14603 ( .B1(n16133), .B2(n16581), .C1(n16134), .C2(n16575), .A(
        n15062), .ZN(n15061) );
  AOI22_X1 U14604 ( .A1(n16569), .A2(n12333), .B1(n16564), .B2(OUT2[56]), .ZN(
        n15062) );
  OAI221_X1 U14605 ( .B1(n7750), .B2(n16635), .C1(n7884), .C2(n16629), .A(
        n15038), .ZN(n15033) );
  AOI22_X1 U14606 ( .A1(n16623), .A2(n13129), .B1(n16617), .B2(n8063), .ZN(
        n15038) );
  OAI221_X1 U14607 ( .B1(n16128), .B2(n16581), .C1(n16129), .C2(n16575), .A(
        n15044), .ZN(n15043) );
  AOI22_X1 U14608 ( .A1(n16569), .A2(n12332), .B1(n16564), .B2(OUT2[57]), .ZN(
        n15044) );
  OAI221_X1 U14609 ( .B1(n7748), .B2(n16635), .C1(n7881), .C2(n16629), .A(
        n15020), .ZN(n15015) );
  AOI22_X1 U14610 ( .A1(n16623), .A2(n13128), .B1(n16617), .B2(n8062), .ZN(
        n15020) );
  OAI221_X1 U14611 ( .B1(n16123), .B2(n16581), .C1(n16124), .C2(n16575), .A(
        n15026), .ZN(n15025) );
  AOI22_X1 U14612 ( .A1(n16569), .A2(n12331), .B1(n16564), .B2(OUT2[58]), .ZN(
        n15026) );
  OAI221_X1 U14613 ( .B1(n7746), .B2(n16635), .C1(n7878), .C2(n16629), .A(
        n15002), .ZN(n14997) );
  AOI22_X1 U14614 ( .A1(n16623), .A2(n13127), .B1(n16617), .B2(n8061), .ZN(
        n15002) );
  OAI221_X1 U14615 ( .B1(n16118), .B2(n16581), .C1(n16119), .C2(n16575), .A(
        n15008), .ZN(n15007) );
  AOI22_X1 U14616 ( .A1(n16569), .A2(n12330), .B1(n16564), .B2(OUT2[59]), .ZN(
        n15008) );
  OAI221_X1 U14617 ( .B1(n7744), .B2(n16636), .C1(n7875), .C2(n16630), .A(
        n14984), .ZN(n14979) );
  AOI22_X1 U14618 ( .A1(n16624), .A2(n13126), .B1(n16618), .B2(n8060), .ZN(
        n14984) );
  OAI221_X1 U14619 ( .B1(n16111), .B2(n16559), .C1(n16112), .C2(n16553), .A(
        n14991), .ZN(n14988) );
  AOI22_X1 U14620 ( .A1(n16542), .A2(n12393), .B1(n16541), .B2(n12265), .ZN(
        n14991) );
  OAI221_X1 U14621 ( .B1(n16113), .B2(n16582), .C1(n16114), .C2(n16576), .A(
        n14990), .ZN(n14989) );
  AOI22_X1 U14622 ( .A1(n16570), .A2(n12329), .B1(n16564), .B2(OUT2[60]), .ZN(
        n14990) );
  OAI221_X1 U14623 ( .B1(n7742), .B2(n16636), .C1(n7872), .C2(n16630), .A(
        n14966), .ZN(n14961) );
  AOI22_X1 U14624 ( .A1(n16624), .A2(n13125), .B1(n16618), .B2(n8059), .ZN(
        n14966) );
  OAI221_X1 U14625 ( .B1(n16106), .B2(n16559), .C1(n16107), .C2(n16553), .A(
        n14973), .ZN(n14970) );
  AOI22_X1 U14626 ( .A1(n16542), .A2(n12392), .B1(n16541), .B2(n12264), .ZN(
        n14973) );
  OAI221_X1 U14627 ( .B1(n16108), .B2(n16582), .C1(n16109), .C2(n16576), .A(
        n14972), .ZN(n14971) );
  AOI22_X1 U14628 ( .A1(n16570), .A2(n12328), .B1(n16564), .B2(OUT2[61]), .ZN(
        n14972) );
  OAI221_X1 U14629 ( .B1(n7740), .B2(n16636), .C1(n7869), .C2(n16630), .A(
        n14948), .ZN(n14943) );
  AOI22_X1 U14630 ( .A1(n16624), .A2(n13124), .B1(n16618), .B2(n8058), .ZN(
        n14948) );
  OAI221_X1 U14631 ( .B1(n16101), .B2(n16559), .C1(n16102), .C2(n16553), .A(
        n14955), .ZN(n14952) );
  AOI22_X1 U14632 ( .A1(n16542), .A2(n12391), .B1(n16541), .B2(n12263), .ZN(
        n14955) );
  OAI221_X1 U14633 ( .B1(n16103), .B2(n16582), .C1(n16104), .C2(n16576), .A(
        n14954), .ZN(n14953) );
  AOI22_X1 U14634 ( .A1(n16570), .A2(n12327), .B1(n16564), .B2(OUT2[62]), .ZN(
        n14954) );
  OAI221_X1 U14635 ( .B1(n7738), .B2(n16636), .C1(n7866), .C2(n16630), .A(
        n14906), .ZN(n14891) );
  AOI22_X1 U14636 ( .A1(n16624), .A2(n13123), .B1(n16618), .B2(n8057), .ZN(
        n14906) );
  OAI221_X1 U14637 ( .B1(n16096), .B2(n16559), .C1(n16097), .C2(n16553), .A(
        n14926), .ZN(n14917) );
  AOI22_X1 U14638 ( .A1(n16542), .A2(n12390), .B1(n16541), .B2(n12262), .ZN(
        n14926) );
  OAI221_X1 U14639 ( .B1(n16098), .B2(n16582), .C1(n16099), .C2(n16576), .A(
        n14921), .ZN(n14918) );
  AOI22_X1 U14640 ( .A1(n16570), .A2(n12326), .B1(n14923), .B2(OUT2[63]), .ZN(
        n14921) );
  OAI221_X1 U14641 ( .B1(n7864), .B2(n16836), .C1(n8055), .C2(n16830), .A(
        n14867), .ZN(n14851) );
  AOI22_X1 U14642 ( .A1(n16824), .A2(n13186), .B1(n16818), .B2(n8120), .ZN(
        n14867) );
  OAI221_X1 U14643 ( .B1(n16413), .B2(n16782), .C1(n16414), .C2(n16776), .A(
        n14873), .ZN(n14872) );
  AOI22_X1 U14644 ( .A1(n16770), .A2(n12389), .B1(n16765), .B2(OUT1[0]), .ZN(
        n14873) );
  OAI221_X1 U14645 ( .B1(n7862), .B2(n16836), .C1(n8052), .C2(n16830), .A(
        n14838), .ZN(n14833) );
  AOI22_X1 U14646 ( .A1(n16824), .A2(n13185), .B1(n16818), .B2(n8119), .ZN(
        n14838) );
  OAI221_X1 U14647 ( .B1(n16408), .B2(n16782), .C1(n16409), .C2(n16776), .A(
        n14844), .ZN(n14843) );
  AOI22_X1 U14648 ( .A1(n16770), .A2(n12388), .B1(n16765), .B2(OUT1[1]), .ZN(
        n14844) );
  OAI221_X1 U14649 ( .B1(n7860), .B2(n16836), .C1(n8049), .C2(n16830), .A(
        n14820), .ZN(n14815) );
  AOI22_X1 U14650 ( .A1(n16824), .A2(n13184), .B1(n16818), .B2(n8118), .ZN(
        n14820) );
  OAI221_X1 U14651 ( .B1(n16403), .B2(n16782), .C1(n16404), .C2(n16776), .A(
        n14826), .ZN(n14825) );
  AOI22_X1 U14652 ( .A1(n16770), .A2(n12387), .B1(n16765), .B2(OUT1[2]), .ZN(
        n14826) );
  OAI221_X1 U14653 ( .B1(n7858), .B2(n16836), .C1(n8046), .C2(n16830), .A(
        n14802), .ZN(n14797) );
  AOI22_X1 U14654 ( .A1(n16824), .A2(n13183), .B1(n16818), .B2(n8117), .ZN(
        n14802) );
  OAI221_X1 U14655 ( .B1(n16398), .B2(n16782), .C1(n16399), .C2(n16776), .A(
        n14808), .ZN(n14807) );
  AOI22_X1 U14656 ( .A1(n16770), .A2(n12386), .B1(n16765), .B2(OUT1[3]), .ZN(
        n14808) );
  OAI221_X1 U14657 ( .B1(n7856), .B2(n16836), .C1(n8043), .C2(n16830), .A(
        n14784), .ZN(n14779) );
  AOI22_X1 U14658 ( .A1(n16824), .A2(n13182), .B1(n16818), .B2(n8116), .ZN(
        n14784) );
  OAI221_X1 U14659 ( .B1(n16393), .B2(n16782), .C1(n16394), .C2(n16776), .A(
        n14790), .ZN(n14789) );
  AOI22_X1 U14660 ( .A1(n16770), .A2(n12385), .B1(n16765), .B2(OUT1[4]), .ZN(
        n14790) );
  OAI221_X1 U14661 ( .B1(n7854), .B2(n16836), .C1(n8040), .C2(n16830), .A(
        n14766), .ZN(n14761) );
  AOI22_X1 U14662 ( .A1(n16824), .A2(n13181), .B1(n16818), .B2(n8115), .ZN(
        n14766) );
  OAI221_X1 U14663 ( .B1(n16388), .B2(n16782), .C1(n16389), .C2(n16776), .A(
        n14772), .ZN(n14771) );
  AOI22_X1 U14664 ( .A1(n16770), .A2(n12384), .B1(n16765), .B2(OUT1[5]), .ZN(
        n14772) );
  OAI221_X1 U14665 ( .B1(n7852), .B2(n16836), .C1(n8037), .C2(n16830), .A(
        n14748), .ZN(n14743) );
  AOI22_X1 U14666 ( .A1(n16824), .A2(n13180), .B1(n16818), .B2(n8114), .ZN(
        n14748) );
  OAI221_X1 U14667 ( .B1(n16383), .B2(n16782), .C1(n16384), .C2(n16776), .A(
        n14754), .ZN(n14753) );
  AOI22_X1 U14668 ( .A1(n16770), .A2(n12383), .B1(n16765), .B2(OUT1[6]), .ZN(
        n14754) );
  OAI221_X1 U14669 ( .B1(n7850), .B2(n16836), .C1(n8034), .C2(n16830), .A(
        n14730), .ZN(n14725) );
  AOI22_X1 U14670 ( .A1(n16824), .A2(n13179), .B1(n16818), .B2(n8113), .ZN(
        n14730) );
  OAI221_X1 U14671 ( .B1(n16378), .B2(n16782), .C1(n16379), .C2(n16776), .A(
        n14736), .ZN(n14735) );
  AOI22_X1 U14672 ( .A1(n16770), .A2(n12382), .B1(n16765), .B2(OUT1[7]), .ZN(
        n14736) );
  OAI221_X1 U14673 ( .B1(n7848), .B2(n16836), .C1(n8031), .C2(n16830), .A(
        n14712), .ZN(n14707) );
  AOI22_X1 U14674 ( .A1(n16824), .A2(n13178), .B1(n16818), .B2(n8112), .ZN(
        n14712) );
  OAI221_X1 U14675 ( .B1(n16373), .B2(n16782), .C1(n16374), .C2(n16776), .A(
        n14718), .ZN(n14717) );
  AOI22_X1 U14676 ( .A1(n16770), .A2(n12381), .B1(n16765), .B2(OUT1[8]), .ZN(
        n14718) );
  OAI221_X1 U14677 ( .B1(n7846), .B2(n16836), .C1(n8028), .C2(n16830), .A(
        n14694), .ZN(n14689) );
  AOI22_X1 U14678 ( .A1(n16824), .A2(n13177), .B1(n16818), .B2(n8111), .ZN(
        n14694) );
  OAI221_X1 U14679 ( .B1(n16368), .B2(n16782), .C1(n16369), .C2(n16776), .A(
        n14700), .ZN(n14699) );
  AOI22_X1 U14680 ( .A1(n16770), .A2(n12380), .B1(n16765), .B2(OUT1[9]), .ZN(
        n14700) );
  OAI221_X1 U14681 ( .B1(n7844), .B2(n16836), .C1(n8025), .C2(n16830), .A(
        n14676), .ZN(n14671) );
  AOI22_X1 U14682 ( .A1(n16824), .A2(n13176), .B1(n16818), .B2(n8110), .ZN(
        n14676) );
  OAI221_X1 U14683 ( .B1(n16363), .B2(n16782), .C1(n16364), .C2(n16776), .A(
        n14682), .ZN(n14681) );
  AOI22_X1 U14684 ( .A1(n16770), .A2(n12379), .B1(n16765), .B2(OUT1[10]), .ZN(
        n14682) );
  OAI221_X1 U14685 ( .B1(n7842), .B2(n16836), .C1(n8022), .C2(n16830), .A(
        n14658), .ZN(n14653) );
  AOI22_X1 U14686 ( .A1(n16824), .A2(n13175), .B1(n16818), .B2(n8109), .ZN(
        n14658) );
  OAI221_X1 U14687 ( .B1(n16358), .B2(n16782), .C1(n16359), .C2(n16776), .A(
        n14664), .ZN(n14663) );
  AOI22_X1 U14688 ( .A1(n16770), .A2(n12378), .B1(n16766), .B2(OUT1[11]), .ZN(
        n14664) );
  OAI221_X1 U14689 ( .B1(n7840), .B2(n16837), .C1(n8019), .C2(n16831), .A(
        n14640), .ZN(n14635) );
  AOI22_X1 U14690 ( .A1(n16825), .A2(n13174), .B1(n16819), .B2(n8108), .ZN(
        n14640) );
  OAI221_X1 U14691 ( .B1(n16353), .B2(n16783), .C1(n16354), .C2(n16777), .A(
        n14646), .ZN(n14645) );
  AOI22_X1 U14692 ( .A1(n16771), .A2(n12377), .B1(n16766), .B2(OUT1[12]), .ZN(
        n14646) );
  OAI221_X1 U14693 ( .B1(n7838), .B2(n16837), .C1(n8016), .C2(n16831), .A(
        n14622), .ZN(n14617) );
  AOI22_X1 U14694 ( .A1(n16825), .A2(n13173), .B1(n16819), .B2(n8107), .ZN(
        n14622) );
  OAI221_X1 U14695 ( .B1(n16348), .B2(n16783), .C1(n16349), .C2(n16777), .A(
        n14628), .ZN(n14627) );
  AOI22_X1 U14696 ( .A1(n16771), .A2(n12376), .B1(n16766), .B2(OUT1[13]), .ZN(
        n14628) );
  OAI221_X1 U14697 ( .B1(n7836), .B2(n16837), .C1(n8013), .C2(n16831), .A(
        n14604), .ZN(n14599) );
  AOI22_X1 U14698 ( .A1(n16825), .A2(n13172), .B1(n16819), .B2(n8106), .ZN(
        n14604) );
  OAI221_X1 U14699 ( .B1(n16343), .B2(n16783), .C1(n16344), .C2(n16777), .A(
        n14610), .ZN(n14609) );
  AOI22_X1 U14700 ( .A1(n16771), .A2(n12375), .B1(n16766), .B2(OUT1[14]), .ZN(
        n14610) );
  OAI221_X1 U14701 ( .B1(n7834), .B2(n16837), .C1(n8010), .C2(n16831), .A(
        n14586), .ZN(n14581) );
  AOI22_X1 U14702 ( .A1(n16825), .A2(n13171), .B1(n16819), .B2(n8105), .ZN(
        n14586) );
  OAI221_X1 U14703 ( .B1(n16338), .B2(n16783), .C1(n16339), .C2(n16777), .A(
        n14592), .ZN(n14591) );
  AOI22_X1 U14704 ( .A1(n16771), .A2(n12374), .B1(n16766), .B2(OUT1[15]), .ZN(
        n14592) );
  OAI221_X1 U14705 ( .B1(n7832), .B2(n16837), .C1(n8007), .C2(n16831), .A(
        n14568), .ZN(n14563) );
  AOI22_X1 U14706 ( .A1(n16825), .A2(n13170), .B1(n16819), .B2(n8104), .ZN(
        n14568) );
  OAI221_X1 U14707 ( .B1(n16333), .B2(n16783), .C1(n16334), .C2(n16777), .A(
        n14574), .ZN(n14573) );
  AOI22_X1 U14708 ( .A1(n16771), .A2(n12373), .B1(n16766), .B2(OUT1[16]), .ZN(
        n14574) );
  OAI221_X1 U14709 ( .B1(n7830), .B2(n16837), .C1(n8004), .C2(n16831), .A(
        n14550), .ZN(n14545) );
  AOI22_X1 U14710 ( .A1(n16825), .A2(n13169), .B1(n16819), .B2(n8103), .ZN(
        n14550) );
  OAI221_X1 U14711 ( .B1(n16328), .B2(n16783), .C1(n16329), .C2(n16777), .A(
        n14556), .ZN(n14555) );
  AOI22_X1 U14712 ( .A1(n16771), .A2(n12372), .B1(n16766), .B2(OUT1[17]), .ZN(
        n14556) );
  OAI221_X1 U14713 ( .B1(n7828), .B2(n16837), .C1(n8001), .C2(n16831), .A(
        n14532), .ZN(n14527) );
  AOI22_X1 U14714 ( .A1(n16825), .A2(n13168), .B1(n16819), .B2(n8102), .ZN(
        n14532) );
  OAI221_X1 U14715 ( .B1(n16323), .B2(n16783), .C1(n16324), .C2(n16777), .A(
        n14538), .ZN(n14537) );
  AOI22_X1 U14716 ( .A1(n16771), .A2(n12371), .B1(n16766), .B2(OUT1[18]), .ZN(
        n14538) );
  OAI221_X1 U14717 ( .B1(n7826), .B2(n16837), .C1(n7998), .C2(n16831), .A(
        n14514), .ZN(n14509) );
  AOI22_X1 U14718 ( .A1(n16825), .A2(n13167), .B1(n16819), .B2(n8101), .ZN(
        n14514) );
  OAI221_X1 U14719 ( .B1(n16318), .B2(n16783), .C1(n16319), .C2(n16777), .A(
        n14520), .ZN(n14519) );
  AOI22_X1 U14720 ( .A1(n16771), .A2(n12370), .B1(n16766), .B2(OUT1[19]), .ZN(
        n14520) );
  OAI221_X1 U14721 ( .B1(n7824), .B2(n16837), .C1(n7995), .C2(n16831), .A(
        n14496), .ZN(n14491) );
  AOI22_X1 U14722 ( .A1(n16825), .A2(n13166), .B1(n16819), .B2(n8100), .ZN(
        n14496) );
  OAI221_X1 U14723 ( .B1(n16313), .B2(n16783), .C1(n16314), .C2(n16777), .A(
        n14502), .ZN(n14501) );
  AOI22_X1 U14724 ( .A1(n16771), .A2(n12369), .B1(n16766), .B2(OUT1[20]), .ZN(
        n14502) );
  OAI221_X1 U14725 ( .B1(n7822), .B2(n16837), .C1(n7992), .C2(n16831), .A(
        n14478), .ZN(n14473) );
  AOI22_X1 U14726 ( .A1(n16825), .A2(n13165), .B1(n16819), .B2(n8099), .ZN(
        n14478) );
  OAI221_X1 U14727 ( .B1(n16308), .B2(n16783), .C1(n16309), .C2(n16777), .A(
        n14484), .ZN(n14483) );
  AOI22_X1 U14728 ( .A1(n16771), .A2(n12368), .B1(n16766), .B2(OUT1[21]), .ZN(
        n14484) );
  OAI221_X1 U14729 ( .B1(n7820), .B2(n16837), .C1(n7989), .C2(n16831), .A(
        n14460), .ZN(n14455) );
  AOI22_X1 U14730 ( .A1(n16825), .A2(n13164), .B1(n16819), .B2(n8098), .ZN(
        n14460) );
  OAI221_X1 U14731 ( .B1(n16303), .B2(n16783), .C1(n16304), .C2(n16777), .A(
        n14466), .ZN(n14465) );
  AOI22_X1 U14732 ( .A1(n16771), .A2(n12367), .B1(n16766), .B2(OUT1[22]), .ZN(
        n14466) );
  OAI221_X1 U14733 ( .B1(n7818), .B2(n16837), .C1(n7986), .C2(n16831), .A(
        n14442), .ZN(n14437) );
  AOI22_X1 U14734 ( .A1(n16825), .A2(n13163), .B1(n16819), .B2(n8097), .ZN(
        n14442) );
  OAI221_X1 U14735 ( .B1(n16298), .B2(n16783), .C1(n16299), .C2(n16777), .A(
        n14448), .ZN(n14447) );
  AOI22_X1 U14736 ( .A1(n16771), .A2(n12366), .B1(n16766), .B2(OUT1[23]), .ZN(
        n14448) );
  OAI221_X1 U14737 ( .B1(n7816), .B2(n16838), .C1(n7983), .C2(n16832), .A(
        n14424), .ZN(n14419) );
  AOI22_X1 U14738 ( .A1(n16826), .A2(n13162), .B1(n16820), .B2(n8096), .ZN(
        n14424) );
  OAI221_X1 U14739 ( .B1(n16293), .B2(n16784), .C1(n16294), .C2(n16778), .A(
        n14430), .ZN(n14429) );
  AOI22_X1 U14740 ( .A1(n16772), .A2(n12365), .B1(n16767), .B2(OUT1[24]), .ZN(
        n14430) );
  OAI221_X1 U14741 ( .B1(n7814), .B2(n16838), .C1(n7980), .C2(n16832), .A(
        n14406), .ZN(n14401) );
  AOI22_X1 U14742 ( .A1(n16826), .A2(n13161), .B1(n16820), .B2(n8095), .ZN(
        n14406) );
  OAI221_X1 U14743 ( .B1(n16288), .B2(n16784), .C1(n16289), .C2(n16778), .A(
        n14412), .ZN(n14411) );
  AOI22_X1 U14744 ( .A1(n16772), .A2(n12364), .B1(n16767), .B2(OUT1[25]), .ZN(
        n14412) );
  OAI221_X1 U14745 ( .B1(n7812), .B2(n16838), .C1(n7977), .C2(n16832), .A(
        n14388), .ZN(n14383) );
  AOI22_X1 U14746 ( .A1(n16826), .A2(n13160), .B1(n16820), .B2(n8094), .ZN(
        n14388) );
  OAI221_X1 U14747 ( .B1(n16283), .B2(n16784), .C1(n16284), .C2(n16778), .A(
        n14394), .ZN(n14393) );
  AOI22_X1 U14748 ( .A1(n16772), .A2(n12363), .B1(n16767), .B2(OUT1[26]), .ZN(
        n14394) );
  OAI221_X1 U14749 ( .B1(n7810), .B2(n16838), .C1(n7974), .C2(n16832), .A(
        n14370), .ZN(n14365) );
  AOI22_X1 U14750 ( .A1(n16826), .A2(n13159), .B1(n16820), .B2(n8093), .ZN(
        n14370) );
  OAI221_X1 U14751 ( .B1(n16278), .B2(n16784), .C1(n16279), .C2(n16778), .A(
        n14376), .ZN(n14375) );
  AOI22_X1 U14752 ( .A1(n16772), .A2(n12362), .B1(n16767), .B2(OUT1[27]), .ZN(
        n14376) );
  OAI221_X1 U14753 ( .B1(n7808), .B2(n16838), .C1(n7971), .C2(n16832), .A(
        n14352), .ZN(n14347) );
  AOI22_X1 U14754 ( .A1(n16826), .A2(n13158), .B1(n16820), .B2(n8092), .ZN(
        n14352) );
  OAI221_X1 U14755 ( .B1(n16273), .B2(n16784), .C1(n16274), .C2(n16778), .A(
        n14358), .ZN(n14357) );
  AOI22_X1 U14756 ( .A1(n16772), .A2(n12361), .B1(n16767), .B2(OUT1[28]), .ZN(
        n14358) );
  OAI221_X1 U14757 ( .B1(n7806), .B2(n16838), .C1(n7968), .C2(n16832), .A(
        n14334), .ZN(n14329) );
  AOI22_X1 U14758 ( .A1(n16826), .A2(n13157), .B1(n16820), .B2(n8091), .ZN(
        n14334) );
  OAI221_X1 U14759 ( .B1(n16268), .B2(n16784), .C1(n16269), .C2(n16778), .A(
        n14340), .ZN(n14339) );
  AOI22_X1 U14760 ( .A1(n16772), .A2(n12360), .B1(n16767), .B2(OUT1[29]), .ZN(
        n14340) );
  OAI221_X1 U14761 ( .B1(n7804), .B2(n16838), .C1(n7965), .C2(n16832), .A(
        n14316), .ZN(n14311) );
  AOI22_X1 U14762 ( .A1(n16826), .A2(n13156), .B1(n16820), .B2(n8090), .ZN(
        n14316) );
  OAI221_X1 U14763 ( .B1(n16263), .B2(n16784), .C1(n16264), .C2(n16778), .A(
        n14322), .ZN(n14321) );
  AOI22_X1 U14764 ( .A1(n16772), .A2(n12359), .B1(n16767), .B2(OUT1[30]), .ZN(
        n14322) );
  OAI221_X1 U14765 ( .B1(n7802), .B2(n16838), .C1(n7962), .C2(n16832), .A(
        n14298), .ZN(n14293) );
  AOI22_X1 U14766 ( .A1(n16826), .A2(n13155), .B1(n16820), .B2(n8089), .ZN(
        n14298) );
  OAI221_X1 U14767 ( .B1(n16258), .B2(n16784), .C1(n16259), .C2(n16778), .A(
        n14304), .ZN(n14303) );
  AOI22_X1 U14768 ( .A1(n16772), .A2(n12358), .B1(n16767), .B2(OUT1[31]), .ZN(
        n14304) );
  OAI221_X1 U14769 ( .B1(n7800), .B2(n16838), .C1(n7959), .C2(n16832), .A(
        n14280), .ZN(n14275) );
  AOI22_X1 U14770 ( .A1(n16826), .A2(n13154), .B1(n16820), .B2(n8088), .ZN(
        n14280) );
  OAI221_X1 U14771 ( .B1(n16253), .B2(n16784), .C1(n16254), .C2(n16778), .A(
        n14286), .ZN(n14285) );
  AOI22_X1 U14772 ( .A1(n16772), .A2(n12357), .B1(n16767), .B2(OUT1[32]), .ZN(
        n14286) );
  OAI221_X1 U14773 ( .B1(n7798), .B2(n16838), .C1(n7956), .C2(n16832), .A(
        n14262), .ZN(n14257) );
  AOI22_X1 U14774 ( .A1(n16826), .A2(n13153), .B1(n16820), .B2(n8087), .ZN(
        n14262) );
  OAI221_X1 U14775 ( .B1(n16248), .B2(n16784), .C1(n16249), .C2(n16778), .A(
        n14268), .ZN(n14267) );
  AOI22_X1 U14776 ( .A1(n16772), .A2(n12356), .B1(n16767), .B2(OUT1[33]), .ZN(
        n14268) );
  OAI221_X1 U14777 ( .B1(n7796), .B2(n16838), .C1(n7953), .C2(n16832), .A(
        n14244), .ZN(n14239) );
  AOI22_X1 U14778 ( .A1(n16826), .A2(n13152), .B1(n16820), .B2(n8086), .ZN(
        n14244) );
  OAI221_X1 U14779 ( .B1(n16243), .B2(n16784), .C1(n16244), .C2(n16778), .A(
        n14250), .ZN(n14249) );
  AOI22_X1 U14780 ( .A1(n16772), .A2(n12355), .B1(n16767), .B2(OUT1[34]), .ZN(
        n14250) );
  OAI221_X1 U14781 ( .B1(n7794), .B2(n16838), .C1(n7950), .C2(n16832), .A(
        n14226), .ZN(n14221) );
  AOI22_X1 U14782 ( .A1(n16826), .A2(n13151), .B1(n16820), .B2(n8085), .ZN(
        n14226) );
  OAI221_X1 U14783 ( .B1(n16238), .B2(n16784), .C1(n16239), .C2(n16778), .A(
        n14232), .ZN(n14231) );
  AOI22_X1 U14784 ( .A1(n16772), .A2(n12354), .B1(n16767), .B2(OUT1[35]), .ZN(
        n14232) );
  OAI221_X1 U14785 ( .B1(n7792), .B2(n16839), .C1(n7947), .C2(n16833), .A(
        n14208), .ZN(n14203) );
  AOI22_X1 U14786 ( .A1(n16827), .A2(n13150), .B1(n16821), .B2(n8084), .ZN(
        n14208) );
  OAI221_X1 U14787 ( .B1(n16233), .B2(n16785), .C1(n16234), .C2(n16779), .A(
        n14214), .ZN(n14213) );
  AOI22_X1 U14788 ( .A1(n16773), .A2(n12353), .B1(n16767), .B2(OUT1[36]), .ZN(
        n14214) );
  OAI221_X1 U14789 ( .B1(n7790), .B2(n16839), .C1(n7944), .C2(n16833), .A(
        n14190), .ZN(n14185) );
  AOI22_X1 U14790 ( .A1(n16827), .A2(n13149), .B1(n16821), .B2(n8083), .ZN(
        n14190) );
  OAI221_X1 U14791 ( .B1(n16228), .B2(n16785), .C1(n16229), .C2(n16779), .A(
        n14196), .ZN(n14195) );
  AOI22_X1 U14792 ( .A1(n16773), .A2(n12352), .B1(n16768), .B2(OUT1[37]), .ZN(
        n14196) );
  OAI221_X1 U14793 ( .B1(n7788), .B2(n16839), .C1(n7941), .C2(n16833), .A(
        n14172), .ZN(n14167) );
  AOI22_X1 U14794 ( .A1(n16827), .A2(n13148), .B1(n16821), .B2(n8082), .ZN(
        n14172) );
  OAI221_X1 U14795 ( .B1(n16223), .B2(n16785), .C1(n16224), .C2(n16779), .A(
        n14178), .ZN(n14177) );
  AOI22_X1 U14796 ( .A1(n16773), .A2(n12351), .B1(n16768), .B2(OUT1[38]), .ZN(
        n14178) );
  OAI221_X1 U14797 ( .B1(n7786), .B2(n16839), .C1(n7938), .C2(n16833), .A(
        n14154), .ZN(n14149) );
  AOI22_X1 U14798 ( .A1(n16827), .A2(n13147), .B1(n16821), .B2(n8081), .ZN(
        n14154) );
  OAI221_X1 U14799 ( .B1(n16218), .B2(n16785), .C1(n16219), .C2(n16779), .A(
        n14160), .ZN(n14159) );
  AOI22_X1 U14800 ( .A1(n16773), .A2(n12350), .B1(n16768), .B2(OUT1[39]), .ZN(
        n14160) );
  OAI221_X1 U14801 ( .B1(n7784), .B2(n16839), .C1(n7935), .C2(n16833), .A(
        n14136), .ZN(n14131) );
  AOI22_X1 U14802 ( .A1(n16827), .A2(n13146), .B1(n16821), .B2(n8080), .ZN(
        n14136) );
  OAI221_X1 U14803 ( .B1(n16213), .B2(n16785), .C1(n16214), .C2(n16779), .A(
        n14142), .ZN(n14141) );
  AOI22_X1 U14804 ( .A1(n16773), .A2(n12349), .B1(n16768), .B2(OUT1[40]), .ZN(
        n14142) );
  OAI221_X1 U14805 ( .B1(n7782), .B2(n16839), .C1(n7932), .C2(n16833), .A(
        n14118), .ZN(n14113) );
  AOI22_X1 U14806 ( .A1(n16827), .A2(n13145), .B1(n16821), .B2(n8079), .ZN(
        n14118) );
  OAI221_X1 U14807 ( .B1(n16208), .B2(n16785), .C1(n16209), .C2(n16779), .A(
        n14124), .ZN(n14123) );
  AOI22_X1 U14808 ( .A1(n16773), .A2(n12348), .B1(n16768), .B2(OUT1[41]), .ZN(
        n14124) );
  OAI221_X1 U14809 ( .B1(n7780), .B2(n16839), .C1(n7929), .C2(n16833), .A(
        n14100), .ZN(n14095) );
  AOI22_X1 U14810 ( .A1(n16827), .A2(n13144), .B1(n16821), .B2(n8078), .ZN(
        n14100) );
  OAI221_X1 U14811 ( .B1(n16203), .B2(n16785), .C1(n16204), .C2(n16779), .A(
        n14106), .ZN(n14105) );
  AOI22_X1 U14812 ( .A1(n16773), .A2(n12347), .B1(n16768), .B2(OUT1[42]), .ZN(
        n14106) );
  OAI221_X1 U14813 ( .B1(n7778), .B2(n16839), .C1(n7926), .C2(n16833), .A(
        n14082), .ZN(n14077) );
  AOI22_X1 U14814 ( .A1(n16827), .A2(n13143), .B1(n16821), .B2(n8077), .ZN(
        n14082) );
  OAI221_X1 U14815 ( .B1(n16198), .B2(n16785), .C1(n16199), .C2(n16779), .A(
        n14088), .ZN(n14087) );
  AOI22_X1 U14816 ( .A1(n16773), .A2(n12346), .B1(n16768), .B2(OUT1[43]), .ZN(
        n14088) );
  OAI221_X1 U14817 ( .B1(n7776), .B2(n16839), .C1(n7923), .C2(n16833), .A(
        n14064), .ZN(n14059) );
  AOI22_X1 U14818 ( .A1(n16827), .A2(n13142), .B1(n16821), .B2(n8076), .ZN(
        n14064) );
  OAI221_X1 U14819 ( .B1(n16193), .B2(n16785), .C1(n16194), .C2(n16779), .A(
        n14070), .ZN(n14069) );
  AOI22_X1 U14820 ( .A1(n16773), .A2(n12345), .B1(n16768), .B2(OUT1[44]), .ZN(
        n14070) );
  OAI221_X1 U14821 ( .B1(n7774), .B2(n16839), .C1(n7920), .C2(n16833), .A(
        n14046), .ZN(n14041) );
  AOI22_X1 U14822 ( .A1(n16827), .A2(n13141), .B1(n16821), .B2(n8075), .ZN(
        n14046) );
  OAI221_X1 U14823 ( .B1(n16188), .B2(n16785), .C1(n16189), .C2(n16779), .A(
        n14052), .ZN(n14051) );
  AOI22_X1 U14824 ( .A1(n16773), .A2(n12344), .B1(n16768), .B2(OUT1[45]), .ZN(
        n14052) );
  OAI221_X1 U14825 ( .B1(n7772), .B2(n16839), .C1(n7917), .C2(n16833), .A(
        n14028), .ZN(n14023) );
  AOI22_X1 U14826 ( .A1(n16827), .A2(n13140), .B1(n16821), .B2(n8074), .ZN(
        n14028) );
  OAI221_X1 U14827 ( .B1(n16183), .B2(n16785), .C1(n16184), .C2(n16779), .A(
        n14034), .ZN(n14033) );
  AOI22_X1 U14828 ( .A1(n16773), .A2(n12343), .B1(n16768), .B2(OUT1[46]), .ZN(
        n14034) );
  OAI221_X1 U14829 ( .B1(n7770), .B2(n16839), .C1(n7914), .C2(n16833), .A(
        n14010), .ZN(n14005) );
  AOI22_X1 U14830 ( .A1(n16827), .A2(n13139), .B1(n16821), .B2(n8073), .ZN(
        n14010) );
  OAI221_X1 U14831 ( .B1(n16178), .B2(n16785), .C1(n16179), .C2(n16779), .A(
        n14016), .ZN(n14015) );
  AOI22_X1 U14832 ( .A1(n16773), .A2(n12342), .B1(n16768), .B2(OUT1[47]), .ZN(
        n14016) );
  OAI221_X1 U14833 ( .B1(n7768), .B2(n16840), .C1(n7911), .C2(n16834), .A(
        n13992), .ZN(n13987) );
  AOI22_X1 U14834 ( .A1(n16828), .A2(n13138), .B1(n16822), .B2(n8072), .ZN(
        n13992) );
  OAI221_X1 U14835 ( .B1(n16173), .B2(n16786), .C1(n16174), .C2(n16780), .A(
        n13998), .ZN(n13997) );
  AOI22_X1 U14836 ( .A1(n16774), .A2(n12341), .B1(n16768), .B2(OUT1[48]), .ZN(
        n13998) );
  OAI221_X1 U14837 ( .B1(n16171), .B2(n16763), .C1(n16172), .C2(n16757), .A(
        n13999), .ZN(n13996) );
  AOI22_X1 U14838 ( .A1(n16751), .A2(n12277), .B1(n16745), .B2(n16467), .ZN(
        n13999) );
  OAI221_X1 U14839 ( .B1(n7766), .B2(n16840), .C1(n7908), .C2(n16834), .A(
        n13974), .ZN(n13969) );
  AOI22_X1 U14840 ( .A1(n16828), .A2(n13137), .B1(n16822), .B2(n8071), .ZN(
        n13974) );
  OAI221_X1 U14841 ( .B1(n16168), .B2(n16786), .C1(n16169), .C2(n16780), .A(
        n13980), .ZN(n13979) );
  AOI22_X1 U14842 ( .A1(n16774), .A2(n12340), .B1(n16768), .B2(OUT1[49]), .ZN(
        n13980) );
  OAI221_X1 U14843 ( .B1(n16166), .B2(n16763), .C1(n16167), .C2(n16757), .A(
        n13981), .ZN(n13978) );
  AOI22_X1 U14844 ( .A1(n16751), .A2(n12276), .B1(n16745), .B2(n16468), .ZN(
        n13981) );
  OAI221_X1 U14845 ( .B1(n7764), .B2(n16840), .C1(n7905), .C2(n16834), .A(
        n13956), .ZN(n13951) );
  AOI22_X1 U14846 ( .A1(n16828), .A2(n13136), .B1(n16822), .B2(n8070), .ZN(
        n13956) );
  OAI221_X1 U14847 ( .B1(n16163), .B2(n16786), .C1(n16164), .C2(n16780), .A(
        n13962), .ZN(n13961) );
  AOI22_X1 U14848 ( .A1(n16774), .A2(n12339), .B1(n16769), .B2(OUT1[50]), .ZN(
        n13962) );
  OAI221_X1 U14849 ( .B1(n16161), .B2(n16763), .C1(n16162), .C2(n16757), .A(
        n13963), .ZN(n13960) );
  AOI22_X1 U14850 ( .A1(n16751), .A2(n12275), .B1(n16745), .B2(n16469), .ZN(
        n13963) );
  OAI221_X1 U14851 ( .B1(n7762), .B2(n16840), .C1(n7902), .C2(n16834), .A(
        n13938), .ZN(n13933) );
  AOI22_X1 U14852 ( .A1(n16828), .A2(n13135), .B1(n16822), .B2(n8069), .ZN(
        n13938) );
  OAI221_X1 U14853 ( .B1(n16158), .B2(n16786), .C1(n16159), .C2(n16780), .A(
        n13944), .ZN(n13943) );
  AOI22_X1 U14854 ( .A1(n16774), .A2(n12338), .B1(n16769), .B2(OUT1[51]), .ZN(
        n13944) );
  OAI221_X1 U14855 ( .B1(n16156), .B2(n16763), .C1(n16157), .C2(n16757), .A(
        n13945), .ZN(n13942) );
  AOI22_X1 U14856 ( .A1(n16751), .A2(n12274), .B1(n16745), .B2(n16470), .ZN(
        n13945) );
  OAI221_X1 U14857 ( .B1(n7760), .B2(n16840), .C1(n7899), .C2(n16834), .A(
        n13920), .ZN(n13915) );
  AOI22_X1 U14858 ( .A1(n16828), .A2(n13134), .B1(n16822), .B2(n8068), .ZN(
        n13920) );
  OAI221_X1 U14859 ( .B1(n16153), .B2(n16786), .C1(n16154), .C2(n16780), .A(
        n13926), .ZN(n13925) );
  AOI22_X1 U14860 ( .A1(n16774), .A2(n12337), .B1(n16769), .B2(OUT1[52]), .ZN(
        n13926) );
  OAI221_X1 U14861 ( .B1(n16151), .B2(n16763), .C1(n16152), .C2(n16757), .A(
        n13927), .ZN(n13924) );
  AOI22_X1 U14862 ( .A1(n16751), .A2(n12273), .B1(n16745), .B2(n16471), .ZN(
        n13927) );
  OAI221_X1 U14863 ( .B1(n7758), .B2(n16840), .C1(n7896), .C2(n16834), .A(
        n13902), .ZN(n13897) );
  AOI22_X1 U14864 ( .A1(n16828), .A2(n13133), .B1(n16822), .B2(n8067), .ZN(
        n13902) );
  OAI221_X1 U14865 ( .B1(n16148), .B2(n16786), .C1(n16149), .C2(n16780), .A(
        n13908), .ZN(n13907) );
  AOI22_X1 U14866 ( .A1(n16774), .A2(n12336), .B1(n16769), .B2(OUT1[53]), .ZN(
        n13908) );
  OAI221_X1 U14867 ( .B1(n16146), .B2(n16763), .C1(n16147), .C2(n16757), .A(
        n13909), .ZN(n13906) );
  AOI22_X1 U14868 ( .A1(n16751), .A2(n12272), .B1(n16745), .B2(n16472), .ZN(
        n13909) );
  OAI221_X1 U14869 ( .B1(n7756), .B2(n16840), .C1(n7893), .C2(n16834), .A(
        n13884), .ZN(n13879) );
  AOI22_X1 U14870 ( .A1(n16828), .A2(n13132), .B1(n16822), .B2(n8066), .ZN(
        n13884) );
  OAI221_X1 U14871 ( .B1(n16143), .B2(n16786), .C1(n16144), .C2(n16780), .A(
        n13890), .ZN(n13889) );
  AOI22_X1 U14872 ( .A1(n16774), .A2(n12335), .B1(n16769), .B2(OUT1[54]), .ZN(
        n13890) );
  OAI221_X1 U14873 ( .B1(n16141), .B2(n16763), .C1(n16142), .C2(n16757), .A(
        n13891), .ZN(n13888) );
  AOI22_X1 U14874 ( .A1(n16751), .A2(n12271), .B1(n16745), .B2(n16473), .ZN(
        n13891) );
  OAI221_X1 U14875 ( .B1(n7754), .B2(n16840), .C1(n7890), .C2(n16834), .A(
        n13866), .ZN(n13861) );
  AOI22_X1 U14876 ( .A1(n16828), .A2(n13131), .B1(n16822), .B2(n8065), .ZN(
        n13866) );
  OAI221_X1 U14877 ( .B1(n16138), .B2(n16786), .C1(n16139), .C2(n16780), .A(
        n13872), .ZN(n13871) );
  AOI22_X1 U14878 ( .A1(n16774), .A2(n12334), .B1(n16769), .B2(OUT1[55]), .ZN(
        n13872) );
  OAI221_X1 U14879 ( .B1(n16136), .B2(n16763), .C1(n16137), .C2(n16757), .A(
        n13873), .ZN(n13870) );
  AOI22_X1 U14880 ( .A1(n16751), .A2(n12270), .B1(n16745), .B2(n16474), .ZN(
        n13873) );
  OAI221_X1 U14881 ( .B1(n7752), .B2(n16840), .C1(n7887), .C2(n16834), .A(
        n13848), .ZN(n13843) );
  AOI22_X1 U14882 ( .A1(n16828), .A2(n13130), .B1(n16822), .B2(n8064), .ZN(
        n13848) );
  OAI221_X1 U14883 ( .B1(n16133), .B2(n16786), .C1(n16134), .C2(n16780), .A(
        n13854), .ZN(n13853) );
  AOI22_X1 U14884 ( .A1(n16774), .A2(n12333), .B1(n16769), .B2(OUT1[56]), .ZN(
        n13854) );
  OAI221_X1 U14885 ( .B1(n16131), .B2(n16763), .C1(n16132), .C2(n16757), .A(
        n13855), .ZN(n13852) );
  AOI22_X1 U14886 ( .A1(n16751), .A2(n12269), .B1(n16745), .B2(n16475), .ZN(
        n13855) );
  OAI221_X1 U14887 ( .B1(n7750), .B2(n16840), .C1(n7884), .C2(n16834), .A(
        n13830), .ZN(n13825) );
  AOI22_X1 U14888 ( .A1(n16828), .A2(n13129), .B1(n16822), .B2(n8063), .ZN(
        n13830) );
  OAI221_X1 U14889 ( .B1(n16128), .B2(n16786), .C1(n16129), .C2(n16780), .A(
        n13836), .ZN(n13835) );
  AOI22_X1 U14890 ( .A1(n16774), .A2(n12332), .B1(n16769), .B2(OUT1[57]), .ZN(
        n13836) );
  OAI221_X1 U14891 ( .B1(n16126), .B2(n16763), .C1(n16127), .C2(n16757), .A(
        n13837), .ZN(n13834) );
  AOI22_X1 U14892 ( .A1(n16751), .A2(n12268), .B1(n16745), .B2(n16476), .ZN(
        n13837) );
  OAI221_X1 U14893 ( .B1(n7748), .B2(n16840), .C1(n7881), .C2(n16834), .A(
        n13812), .ZN(n13807) );
  AOI22_X1 U14894 ( .A1(n16828), .A2(n13128), .B1(n16822), .B2(n8062), .ZN(
        n13812) );
  OAI221_X1 U14895 ( .B1(n16123), .B2(n16786), .C1(n16124), .C2(n16780), .A(
        n13818), .ZN(n13817) );
  AOI22_X1 U14896 ( .A1(n16774), .A2(n12331), .B1(n16769), .B2(OUT1[58]), .ZN(
        n13818) );
  OAI221_X1 U14897 ( .B1(n16121), .B2(n16763), .C1(n16122), .C2(n16757), .A(
        n13819), .ZN(n13816) );
  AOI22_X1 U14898 ( .A1(n16751), .A2(n12267), .B1(n16745), .B2(n16477), .ZN(
        n13819) );
  OAI221_X1 U14899 ( .B1(n7746), .B2(n16840), .C1(n7878), .C2(n16834), .A(
        n13794), .ZN(n13789) );
  AOI22_X1 U14900 ( .A1(n16828), .A2(n13127), .B1(n16822), .B2(n8061), .ZN(
        n13794) );
  OAI221_X1 U14901 ( .B1(n16118), .B2(n16786), .C1(n16119), .C2(n16780), .A(
        n13800), .ZN(n13799) );
  AOI22_X1 U14902 ( .A1(n16774), .A2(n12330), .B1(n16769), .B2(OUT1[59]), .ZN(
        n13800) );
  OAI221_X1 U14903 ( .B1(n16116), .B2(n16763), .C1(n16117), .C2(n16757), .A(
        n13801), .ZN(n13798) );
  AOI22_X1 U14904 ( .A1(n16751), .A2(n12266), .B1(n16745), .B2(n16478), .ZN(
        n13801) );
  OAI221_X1 U14905 ( .B1(n7744), .B2(n16841), .C1(n7875), .C2(n16835), .A(
        n13776), .ZN(n13771) );
  AOI22_X1 U14906 ( .A1(n16829), .A2(n13126), .B1(n16823), .B2(n8060), .ZN(
        n13776) );
  OAI221_X1 U14907 ( .B1(n16113), .B2(n16787), .C1(n16114), .C2(n16781), .A(
        n13782), .ZN(n13781) );
  AOI22_X1 U14908 ( .A1(n16775), .A2(n12329), .B1(n16769), .B2(OUT1[60]), .ZN(
        n13782) );
  OAI221_X1 U14909 ( .B1(n16111), .B2(n16764), .C1(n16112), .C2(n16758), .A(
        n13783), .ZN(n13780) );
  AOI22_X1 U14910 ( .A1(n16752), .A2(n12265), .B1(n16746), .B2(n16416), .ZN(
        n13783) );
  OAI221_X1 U14911 ( .B1(n7742), .B2(n16841), .C1(n7872), .C2(n16835), .A(
        n13758), .ZN(n13753) );
  AOI22_X1 U14912 ( .A1(n16829), .A2(n13125), .B1(n16823), .B2(n8059), .ZN(
        n13758) );
  OAI221_X1 U14913 ( .B1(n16108), .B2(n16787), .C1(n16109), .C2(n16781), .A(
        n13764), .ZN(n13763) );
  AOI22_X1 U14914 ( .A1(n16775), .A2(n12328), .B1(n16769), .B2(OUT1[61]), .ZN(
        n13764) );
  OAI221_X1 U14915 ( .B1(n16106), .B2(n16764), .C1(n16107), .C2(n16758), .A(
        n13765), .ZN(n13762) );
  AOI22_X1 U14916 ( .A1(n16752), .A2(n12264), .B1(n16746), .B2(n16417), .ZN(
        n13765) );
  OAI221_X1 U14917 ( .B1(n7740), .B2(n16841), .C1(n7869), .C2(n16835), .A(
        n13740), .ZN(n13735) );
  AOI22_X1 U14918 ( .A1(n16829), .A2(n13124), .B1(n16823), .B2(n8058), .ZN(
        n13740) );
  OAI221_X1 U14919 ( .B1(n16103), .B2(n16787), .C1(n16104), .C2(n16781), .A(
        n13746), .ZN(n13745) );
  AOI22_X1 U14920 ( .A1(n16775), .A2(n12327), .B1(n16769), .B2(OUT1[62]), .ZN(
        n13746) );
  OAI221_X1 U14921 ( .B1(n16101), .B2(n16764), .C1(n16102), .C2(n16758), .A(
        n13747), .ZN(n13744) );
  AOI22_X1 U14922 ( .A1(n16752), .A2(n12263), .B1(n16746), .B2(n16418), .ZN(
        n13747) );
  OAI221_X1 U14923 ( .B1(n7738), .B2(n16841), .C1(n7866), .C2(n16835), .A(
        n13698), .ZN(n13683) );
  AOI22_X1 U14924 ( .A1(n16829), .A2(n13123), .B1(n16823), .B2(n8057), .ZN(
        n13698) );
  OAI221_X1 U14925 ( .B1(n16098), .B2(n16787), .C1(n16099), .C2(n16781), .A(
        n13713), .ZN(n13710) );
  AOI22_X1 U14926 ( .A1(n16775), .A2(n12326), .B1(n13715), .B2(OUT1[63]), .ZN(
        n13713) );
  OAI221_X1 U14927 ( .B1(n16096), .B2(n16764), .C1(n16097), .C2(n16758), .A(
        n13718), .ZN(n13709) );
  AOI22_X1 U14928 ( .A1(n16752), .A2(n12262), .B1(n16746), .B2(n16419), .ZN(
        n13718) );
  OAI22_X1 U14929 ( .A1(n16965), .A2(n17480), .B1(n16959), .B2(n13354), .ZN(
        n5284) );
  OAI22_X1 U14930 ( .A1(n16966), .A2(n17482), .B1(n16960), .B2(n13353), .ZN(
        n5285) );
  OAI22_X1 U14931 ( .A1(n16966), .A2(n17484), .B1(n16958), .B2(n13352), .ZN(
        n5286) );
  OAI22_X1 U14932 ( .A1(n16966), .A2(n17486), .B1(n16959), .B2(n13351), .ZN(
        n5287) );
  OAI22_X1 U14933 ( .A1(n16966), .A2(n17488), .B1(n16960), .B2(n13350), .ZN(
        n5288) );
  OAI22_X1 U14934 ( .A1(n16966), .A2(n17490), .B1(n16958), .B2(n13349), .ZN(
        n5289) );
  OAI22_X1 U14935 ( .A1(n16967), .A2(n17492), .B1(n16959), .B2(n13348), .ZN(
        n5290) );
  OAI22_X1 U14936 ( .A1(n16967), .A2(n17494), .B1(n16960), .B2(n13347), .ZN(
        n5291) );
  OAI22_X1 U14937 ( .A1(n16967), .A2(n17496), .B1(n16958), .B2(n13346), .ZN(
        n5292) );
  OAI22_X1 U14938 ( .A1(n16967), .A2(n17498), .B1(n16959), .B2(n13345), .ZN(
        n5293) );
  OAI22_X1 U14939 ( .A1(n16967), .A2(n17500), .B1(n16960), .B2(n13344), .ZN(
        n5294) );
  OAI22_X1 U14940 ( .A1(n16968), .A2(n17502), .B1(n16958), .B2(n13343), .ZN(
        n5295) );
  OAI22_X1 U14941 ( .A1(n16968), .A2(n17504), .B1(n13675), .B2(n13342), .ZN(
        n5296) );
  OAI22_X1 U14942 ( .A1(n16968), .A2(n17506), .B1(n16958), .B2(n13341), .ZN(
        n5297) );
  OAI22_X1 U14943 ( .A1(n16968), .A2(n17508), .B1(n13675), .B2(n13340), .ZN(
        n5298) );
  OAI22_X1 U14944 ( .A1(n16968), .A2(n17510), .B1(n16958), .B2(n13339), .ZN(
        n5299) );
  OAI22_X1 U14945 ( .A1(n16969), .A2(n17512), .B1(n13675), .B2(n13338), .ZN(
        n5300) );
  OAI22_X1 U14946 ( .A1(n16969), .A2(n17514), .B1(n16958), .B2(n13337), .ZN(
        n5301) );
  OAI22_X1 U14947 ( .A1(n16969), .A2(n17516), .B1(n16959), .B2(n13336), .ZN(
        n5302) );
  OAI22_X1 U14948 ( .A1(n16969), .A2(n17518), .B1(n16960), .B2(n13335), .ZN(
        n5303) );
  OAI22_X1 U14949 ( .A1(n16969), .A2(n17520), .B1(n16958), .B2(n13334), .ZN(
        n5304) );
  OAI22_X1 U14950 ( .A1(n16970), .A2(n17522), .B1(n16958), .B2(n13333), .ZN(
        n5305) );
  OAI22_X1 U14951 ( .A1(n16970), .A2(n17524), .B1(n16959), .B2(n13332), .ZN(
        n5306) );
  OAI22_X1 U14952 ( .A1(n16970), .A2(n17526), .B1(n16960), .B2(n13331), .ZN(
        n5307) );
  OAI22_X1 U14953 ( .A1(n16970), .A2(n17528), .B1(n16958), .B2(n13330), .ZN(
        n5308) );
  OAI22_X1 U14954 ( .A1(n16970), .A2(n17530), .B1(n16958), .B2(n13329), .ZN(
        n5309) );
  OAI22_X1 U14955 ( .A1(n16971), .A2(n17532), .B1(n13675), .B2(n13328), .ZN(
        n5310) );
  OAI22_X1 U14956 ( .A1(n16971), .A2(n17534), .B1(n16958), .B2(n13327), .ZN(
        n5311) );
  OAI22_X1 U14957 ( .A1(n16971), .A2(n17536), .B1(n13675), .B2(n13326), .ZN(
        n5312) );
  OAI22_X1 U14958 ( .A1(n16971), .A2(n17538), .B1(n16958), .B2(n13325), .ZN(
        n5313) );
  OAI22_X1 U14959 ( .A1(n16971), .A2(n17540), .B1(n13675), .B2(n13324), .ZN(
        n5314) );
  OAI22_X1 U14960 ( .A1(n16972), .A2(n17542), .B1(n16958), .B2(n13323), .ZN(
        n5315) );
  OAI22_X1 U14961 ( .A1(n16972), .A2(n17544), .B1(n13675), .B2(n13322), .ZN(
        n5316) );
  OAI22_X1 U14962 ( .A1(n16972), .A2(n17546), .B1(n16958), .B2(n13321), .ZN(
        n5317) );
  OAI22_X1 U14963 ( .A1(n16972), .A2(n17548), .B1(n13675), .B2(n13320), .ZN(
        n5318) );
  OAI22_X1 U14964 ( .A1(n16972), .A2(n17550), .B1(n16958), .B2(n13319), .ZN(
        n5319) );
  OAI22_X1 U14965 ( .A1(n16982), .A2(n17480), .B1(n16976), .B2(n13290), .ZN(
        n5348) );
  OAI22_X1 U14966 ( .A1(n16983), .A2(n17482), .B1(n16977), .B2(n13289), .ZN(
        n5349) );
  OAI22_X1 U14967 ( .A1(n16983), .A2(n17484), .B1(n16975), .B2(n13288), .ZN(
        n5350) );
  OAI22_X1 U14968 ( .A1(n16983), .A2(n17486), .B1(n16976), .B2(n13287), .ZN(
        n5351) );
  OAI22_X1 U14969 ( .A1(n16983), .A2(n17488), .B1(n16977), .B2(n13286), .ZN(
        n5352) );
  OAI22_X1 U14970 ( .A1(n16983), .A2(n17490), .B1(n16975), .B2(n13285), .ZN(
        n5353) );
  OAI22_X1 U14971 ( .A1(n16984), .A2(n17492), .B1(n16976), .B2(n13284), .ZN(
        n5354) );
  OAI22_X1 U14972 ( .A1(n16984), .A2(n17494), .B1(n16977), .B2(n13283), .ZN(
        n5355) );
  OAI22_X1 U14973 ( .A1(n16984), .A2(n17496), .B1(n16975), .B2(n13282), .ZN(
        n5356) );
  OAI22_X1 U14974 ( .A1(n16984), .A2(n17498), .B1(n16976), .B2(n13281), .ZN(
        n5357) );
  OAI22_X1 U14975 ( .A1(n16984), .A2(n17500), .B1(n16977), .B2(n13280), .ZN(
        n5358) );
  OAI22_X1 U14976 ( .A1(n16985), .A2(n17502), .B1(n16975), .B2(n13279), .ZN(
        n5359) );
  OAI22_X1 U14977 ( .A1(n16985), .A2(n17504), .B1(n13674), .B2(n13278), .ZN(
        n5360) );
  OAI22_X1 U14978 ( .A1(n16985), .A2(n17506), .B1(n16975), .B2(n13277), .ZN(
        n5361) );
  OAI22_X1 U14979 ( .A1(n16985), .A2(n17508), .B1(n13674), .B2(n13276), .ZN(
        n5362) );
  OAI22_X1 U14980 ( .A1(n16985), .A2(n17510), .B1(n16975), .B2(n13275), .ZN(
        n5363) );
  OAI22_X1 U14981 ( .A1(n16986), .A2(n17512), .B1(n13674), .B2(n13274), .ZN(
        n5364) );
  OAI22_X1 U14982 ( .A1(n16986), .A2(n17514), .B1(n16975), .B2(n13273), .ZN(
        n5365) );
  OAI22_X1 U14983 ( .A1(n16986), .A2(n17516), .B1(n16976), .B2(n13272), .ZN(
        n5366) );
  OAI22_X1 U14984 ( .A1(n16986), .A2(n17518), .B1(n16977), .B2(n13271), .ZN(
        n5367) );
  OAI22_X1 U14985 ( .A1(n16986), .A2(n17520), .B1(n16975), .B2(n13270), .ZN(
        n5368) );
  OAI22_X1 U14986 ( .A1(n16987), .A2(n17522), .B1(n16975), .B2(n13269), .ZN(
        n5369) );
  OAI22_X1 U14987 ( .A1(n16987), .A2(n17524), .B1(n16976), .B2(n13268), .ZN(
        n5370) );
  OAI22_X1 U14988 ( .A1(n16987), .A2(n17526), .B1(n16977), .B2(n13267), .ZN(
        n5371) );
  OAI22_X1 U14989 ( .A1(n16987), .A2(n17528), .B1(n16975), .B2(n13266), .ZN(
        n5372) );
  OAI22_X1 U14990 ( .A1(n16987), .A2(n17530), .B1(n16975), .B2(n13265), .ZN(
        n5373) );
  OAI22_X1 U14991 ( .A1(n16988), .A2(n17532), .B1(n13674), .B2(n13264), .ZN(
        n5374) );
  OAI22_X1 U14992 ( .A1(n16988), .A2(n17534), .B1(n16975), .B2(n13263), .ZN(
        n5375) );
  OAI22_X1 U14993 ( .A1(n16988), .A2(n17536), .B1(n13674), .B2(n13262), .ZN(
        n5376) );
  OAI22_X1 U14994 ( .A1(n16988), .A2(n17538), .B1(n16975), .B2(n13261), .ZN(
        n5377) );
  OAI22_X1 U14995 ( .A1(n16988), .A2(n17540), .B1(n13674), .B2(n13260), .ZN(
        n5378) );
  OAI22_X1 U14996 ( .A1(n16989), .A2(n17542), .B1(n16975), .B2(n13259), .ZN(
        n5379) );
  OAI22_X1 U14997 ( .A1(n16989), .A2(n17544), .B1(n13674), .B2(n13258), .ZN(
        n5380) );
  OAI22_X1 U14998 ( .A1(n16989), .A2(n17546), .B1(n16975), .B2(n13257), .ZN(
        n5381) );
  OAI22_X1 U14999 ( .A1(n16989), .A2(n17548), .B1(n13674), .B2(n13256), .ZN(
        n5382) );
  OAI22_X1 U15000 ( .A1(n16989), .A2(n17550), .B1(n16975), .B2(n13255), .ZN(
        n5383) );
  OAI22_X1 U15001 ( .A1(n17084), .A2(n17480), .B1(n17078), .B2(n12970), .ZN(
        n5732) );
  OAI22_X1 U15002 ( .A1(n17085), .A2(n17482), .B1(n17079), .B2(n12969), .ZN(
        n5733) );
  OAI22_X1 U15003 ( .A1(n17085), .A2(n17484), .B1(n17077), .B2(n12968), .ZN(
        n5734) );
  OAI22_X1 U15004 ( .A1(n17085), .A2(n17486), .B1(n17078), .B2(n12967), .ZN(
        n5735) );
  OAI22_X1 U15005 ( .A1(n17085), .A2(n17488), .B1(n17079), .B2(n12966), .ZN(
        n5736) );
  OAI22_X1 U15006 ( .A1(n17085), .A2(n17490), .B1(n17077), .B2(n12965), .ZN(
        n5737) );
  OAI22_X1 U15007 ( .A1(n17086), .A2(n17492), .B1(n17078), .B2(n12964), .ZN(
        n5738) );
  OAI22_X1 U15008 ( .A1(n17086), .A2(n17494), .B1(n17079), .B2(n12963), .ZN(
        n5739) );
  OAI22_X1 U15009 ( .A1(n17086), .A2(n17496), .B1(n17077), .B2(n12962), .ZN(
        n5740) );
  OAI22_X1 U15010 ( .A1(n17086), .A2(n17498), .B1(n17078), .B2(n12961), .ZN(
        n5741) );
  OAI22_X1 U15011 ( .A1(n17086), .A2(n17500), .B1(n17079), .B2(n12960), .ZN(
        n5742) );
  OAI22_X1 U15012 ( .A1(n17087), .A2(n17502), .B1(n17077), .B2(n12959), .ZN(
        n5743) );
  OAI22_X1 U15013 ( .A1(n17087), .A2(n17504), .B1(n13667), .B2(n12958), .ZN(
        n5744) );
  OAI22_X1 U15014 ( .A1(n17087), .A2(n17506), .B1(n17077), .B2(n12957), .ZN(
        n5745) );
  OAI22_X1 U15015 ( .A1(n17087), .A2(n17508), .B1(n13667), .B2(n12956), .ZN(
        n5746) );
  OAI22_X1 U15016 ( .A1(n17087), .A2(n17510), .B1(n17077), .B2(n12955), .ZN(
        n5747) );
  OAI22_X1 U15017 ( .A1(n17088), .A2(n17512), .B1(n13667), .B2(n12954), .ZN(
        n5748) );
  OAI22_X1 U15018 ( .A1(n17088), .A2(n17514), .B1(n17077), .B2(n12953), .ZN(
        n5749) );
  OAI22_X1 U15019 ( .A1(n17088), .A2(n17516), .B1(n17078), .B2(n12952), .ZN(
        n5750) );
  OAI22_X1 U15020 ( .A1(n17088), .A2(n17518), .B1(n17079), .B2(n12951), .ZN(
        n5751) );
  OAI22_X1 U15021 ( .A1(n17088), .A2(n17520), .B1(n17077), .B2(n12950), .ZN(
        n5752) );
  OAI22_X1 U15022 ( .A1(n17089), .A2(n17522), .B1(n17077), .B2(n12949), .ZN(
        n5753) );
  OAI22_X1 U15023 ( .A1(n17089), .A2(n17524), .B1(n17078), .B2(n12948), .ZN(
        n5754) );
  OAI22_X1 U15024 ( .A1(n17089), .A2(n17526), .B1(n17079), .B2(n12947), .ZN(
        n5755) );
  OAI22_X1 U15025 ( .A1(n17089), .A2(n17528), .B1(n17077), .B2(n12946), .ZN(
        n5756) );
  OAI22_X1 U15026 ( .A1(n17089), .A2(n17530), .B1(n17077), .B2(n12945), .ZN(
        n5757) );
  OAI22_X1 U15027 ( .A1(n17090), .A2(n17532), .B1(n13667), .B2(n12944), .ZN(
        n5758) );
  OAI22_X1 U15028 ( .A1(n17090), .A2(n17534), .B1(n17077), .B2(n12943), .ZN(
        n5759) );
  OAI22_X1 U15029 ( .A1(n17090), .A2(n17536), .B1(n13667), .B2(n12942), .ZN(
        n5760) );
  OAI22_X1 U15030 ( .A1(n17090), .A2(n17538), .B1(n17077), .B2(n12941), .ZN(
        n5761) );
  OAI22_X1 U15031 ( .A1(n17090), .A2(n17540), .B1(n13667), .B2(n12940), .ZN(
        n5762) );
  OAI22_X1 U15032 ( .A1(n17091), .A2(n17542), .B1(n17077), .B2(n12939), .ZN(
        n5763) );
  OAI22_X1 U15033 ( .A1(n17091), .A2(n17544), .B1(n13667), .B2(n12938), .ZN(
        n5764) );
  OAI22_X1 U15034 ( .A1(n17091), .A2(n17546), .B1(n17077), .B2(n12937), .ZN(
        n5765) );
  OAI22_X1 U15035 ( .A1(n17091), .A2(n17548), .B1(n13667), .B2(n12936), .ZN(
        n5766) );
  OAI22_X1 U15036 ( .A1(n17091), .A2(n17550), .B1(n17077), .B2(n12935), .ZN(
        n5767) );
  OAI22_X1 U15037 ( .A1(n17135), .A2(n17481), .B1(n17129), .B2(n12906), .ZN(
        n5924) );
  OAI22_X1 U15038 ( .A1(n17136), .A2(n17483), .B1(n17130), .B2(n12905), .ZN(
        n5925) );
  OAI22_X1 U15039 ( .A1(n17136), .A2(n17485), .B1(n17128), .B2(n12904), .ZN(
        n5926) );
  OAI22_X1 U15040 ( .A1(n17136), .A2(n17487), .B1(n17129), .B2(n12903), .ZN(
        n5927) );
  OAI22_X1 U15041 ( .A1(n17136), .A2(n17489), .B1(n17130), .B2(n12902), .ZN(
        n5928) );
  OAI22_X1 U15042 ( .A1(n17136), .A2(n17491), .B1(n17128), .B2(n12901), .ZN(
        n5929) );
  OAI22_X1 U15043 ( .A1(n17137), .A2(n17493), .B1(n17129), .B2(n12900), .ZN(
        n5930) );
  OAI22_X1 U15044 ( .A1(n17137), .A2(n17495), .B1(n17130), .B2(n12899), .ZN(
        n5931) );
  OAI22_X1 U15045 ( .A1(n17137), .A2(n17497), .B1(n17128), .B2(n12898), .ZN(
        n5932) );
  OAI22_X1 U15046 ( .A1(n17137), .A2(n17499), .B1(n17129), .B2(n12897), .ZN(
        n5933) );
  OAI22_X1 U15047 ( .A1(n17137), .A2(n17501), .B1(n17130), .B2(n12896), .ZN(
        n5934) );
  OAI22_X1 U15048 ( .A1(n17138), .A2(n17503), .B1(n17128), .B2(n12895), .ZN(
        n5935) );
  OAI22_X1 U15049 ( .A1(n17138), .A2(n17505), .B1(n13664), .B2(n12894), .ZN(
        n5936) );
  OAI22_X1 U15050 ( .A1(n17138), .A2(n17507), .B1(n17128), .B2(n12893), .ZN(
        n5937) );
  OAI22_X1 U15051 ( .A1(n17138), .A2(n17509), .B1(n13664), .B2(n12892), .ZN(
        n5938) );
  OAI22_X1 U15052 ( .A1(n17138), .A2(n17511), .B1(n17128), .B2(n12891), .ZN(
        n5939) );
  OAI22_X1 U15053 ( .A1(n17139), .A2(n17513), .B1(n13664), .B2(n12890), .ZN(
        n5940) );
  OAI22_X1 U15054 ( .A1(n17139), .A2(n17515), .B1(n17128), .B2(n12889), .ZN(
        n5941) );
  OAI22_X1 U15055 ( .A1(n17139), .A2(n17517), .B1(n17129), .B2(n12888), .ZN(
        n5942) );
  OAI22_X1 U15056 ( .A1(n17139), .A2(n17519), .B1(n17130), .B2(n12887), .ZN(
        n5943) );
  OAI22_X1 U15057 ( .A1(n17139), .A2(n17521), .B1(n17128), .B2(n12886), .ZN(
        n5944) );
  OAI22_X1 U15058 ( .A1(n17140), .A2(n17523), .B1(n17128), .B2(n12885), .ZN(
        n5945) );
  OAI22_X1 U15059 ( .A1(n17140), .A2(n17525), .B1(n17129), .B2(n12884), .ZN(
        n5946) );
  OAI22_X1 U15060 ( .A1(n17140), .A2(n17527), .B1(n17130), .B2(n12883), .ZN(
        n5947) );
  OAI22_X1 U15061 ( .A1(n17140), .A2(n17529), .B1(n17128), .B2(n12882), .ZN(
        n5948) );
  OAI22_X1 U15062 ( .A1(n17140), .A2(n17531), .B1(n17128), .B2(n12881), .ZN(
        n5949) );
  OAI22_X1 U15063 ( .A1(n17141), .A2(n17533), .B1(n13664), .B2(n12880), .ZN(
        n5950) );
  OAI22_X1 U15064 ( .A1(n17141), .A2(n17535), .B1(n17128), .B2(n12879), .ZN(
        n5951) );
  OAI22_X1 U15065 ( .A1(n17141), .A2(n17537), .B1(n13664), .B2(n12878), .ZN(
        n5952) );
  OAI22_X1 U15066 ( .A1(n17141), .A2(n17539), .B1(n17128), .B2(n12877), .ZN(
        n5953) );
  OAI22_X1 U15067 ( .A1(n17141), .A2(n17541), .B1(n13664), .B2(n12876), .ZN(
        n5954) );
  OAI22_X1 U15068 ( .A1(n17142), .A2(n17543), .B1(n17128), .B2(n12875), .ZN(
        n5955) );
  OAI22_X1 U15069 ( .A1(n17142), .A2(n17545), .B1(n13664), .B2(n12874), .ZN(
        n5956) );
  OAI22_X1 U15070 ( .A1(n17142), .A2(n17547), .B1(n17128), .B2(n12873), .ZN(
        n5957) );
  OAI22_X1 U15071 ( .A1(n17142), .A2(n17549), .B1(n13664), .B2(n12872), .ZN(
        n5958) );
  OAI22_X1 U15072 ( .A1(n17142), .A2(n17551), .B1(n17128), .B2(n12871), .ZN(
        n5959) );
  OAI22_X1 U15073 ( .A1(n17152), .A2(n17481), .B1(n17146), .B2(n12842), .ZN(
        n5988) );
  OAI22_X1 U15074 ( .A1(n17153), .A2(n17483), .B1(n17147), .B2(n12841), .ZN(
        n5989) );
  OAI22_X1 U15075 ( .A1(n17153), .A2(n17485), .B1(n17145), .B2(n12840), .ZN(
        n5990) );
  OAI22_X1 U15076 ( .A1(n17153), .A2(n17487), .B1(n17146), .B2(n12839), .ZN(
        n5991) );
  OAI22_X1 U15077 ( .A1(n17153), .A2(n17489), .B1(n17147), .B2(n12838), .ZN(
        n5992) );
  OAI22_X1 U15078 ( .A1(n17153), .A2(n17491), .B1(n17145), .B2(n12837), .ZN(
        n5993) );
  OAI22_X1 U15079 ( .A1(n17154), .A2(n17493), .B1(n17146), .B2(n12836), .ZN(
        n5994) );
  OAI22_X1 U15080 ( .A1(n17154), .A2(n17495), .B1(n17147), .B2(n12835), .ZN(
        n5995) );
  OAI22_X1 U15081 ( .A1(n17154), .A2(n17497), .B1(n17145), .B2(n12834), .ZN(
        n5996) );
  OAI22_X1 U15082 ( .A1(n17154), .A2(n17499), .B1(n17146), .B2(n12833), .ZN(
        n5997) );
  OAI22_X1 U15083 ( .A1(n17154), .A2(n17501), .B1(n17147), .B2(n12832), .ZN(
        n5998) );
  OAI22_X1 U15084 ( .A1(n17155), .A2(n17503), .B1(n17145), .B2(n12831), .ZN(
        n5999) );
  OAI22_X1 U15085 ( .A1(n17155), .A2(n17505), .B1(n13662), .B2(n12830), .ZN(
        n6000) );
  OAI22_X1 U15086 ( .A1(n17155), .A2(n17507), .B1(n17145), .B2(n12829), .ZN(
        n6001) );
  OAI22_X1 U15087 ( .A1(n17155), .A2(n17509), .B1(n13662), .B2(n12828), .ZN(
        n6002) );
  OAI22_X1 U15088 ( .A1(n17155), .A2(n17511), .B1(n17145), .B2(n12827), .ZN(
        n6003) );
  OAI22_X1 U15089 ( .A1(n17156), .A2(n17513), .B1(n13662), .B2(n12826), .ZN(
        n6004) );
  OAI22_X1 U15090 ( .A1(n17156), .A2(n17515), .B1(n17145), .B2(n12825), .ZN(
        n6005) );
  OAI22_X1 U15091 ( .A1(n17156), .A2(n17517), .B1(n17146), .B2(n12824), .ZN(
        n6006) );
  OAI22_X1 U15092 ( .A1(n17156), .A2(n17519), .B1(n17147), .B2(n12823), .ZN(
        n6007) );
  OAI22_X1 U15093 ( .A1(n17156), .A2(n17521), .B1(n17145), .B2(n12822), .ZN(
        n6008) );
  OAI22_X1 U15094 ( .A1(n17157), .A2(n17523), .B1(n17145), .B2(n12821), .ZN(
        n6009) );
  OAI22_X1 U15095 ( .A1(n17157), .A2(n17525), .B1(n17146), .B2(n12820), .ZN(
        n6010) );
  OAI22_X1 U15096 ( .A1(n17157), .A2(n17527), .B1(n17147), .B2(n12819), .ZN(
        n6011) );
  OAI22_X1 U15097 ( .A1(n17157), .A2(n17529), .B1(n17145), .B2(n12818), .ZN(
        n6012) );
  OAI22_X1 U15098 ( .A1(n17157), .A2(n17531), .B1(n17145), .B2(n12817), .ZN(
        n6013) );
  OAI22_X1 U15099 ( .A1(n17158), .A2(n17533), .B1(n13662), .B2(n12816), .ZN(
        n6014) );
  OAI22_X1 U15100 ( .A1(n17158), .A2(n17535), .B1(n17145), .B2(n12815), .ZN(
        n6015) );
  OAI22_X1 U15101 ( .A1(n17158), .A2(n17537), .B1(n13662), .B2(n12814), .ZN(
        n6016) );
  OAI22_X1 U15102 ( .A1(n17158), .A2(n17539), .B1(n17145), .B2(n12813), .ZN(
        n6017) );
  OAI22_X1 U15103 ( .A1(n17158), .A2(n17541), .B1(n13662), .B2(n12812), .ZN(
        n6018) );
  OAI22_X1 U15104 ( .A1(n17159), .A2(n17543), .B1(n17145), .B2(n12811), .ZN(
        n6019) );
  OAI22_X1 U15105 ( .A1(n17159), .A2(n17545), .B1(n13662), .B2(n12810), .ZN(
        n6020) );
  OAI22_X1 U15106 ( .A1(n17159), .A2(n17547), .B1(n17145), .B2(n12809), .ZN(
        n6021) );
  OAI22_X1 U15107 ( .A1(n17159), .A2(n17549), .B1(n13662), .B2(n12808), .ZN(
        n6022) );
  OAI22_X1 U15108 ( .A1(n17159), .A2(n17551), .B1(n17145), .B2(n12807), .ZN(
        n6023) );
  OAI22_X1 U15109 ( .A1(n17272), .A2(n17481), .B1(n17266), .B2(n12557), .ZN(
        n6436) );
  OAI22_X1 U15110 ( .A1(n17273), .A2(n17483), .B1(n17267), .B2(n12556), .ZN(
        n6437) );
  OAI22_X1 U15111 ( .A1(n17273), .A2(n17485), .B1(n17265), .B2(n12555), .ZN(
        n6438) );
  OAI22_X1 U15112 ( .A1(n17273), .A2(n17487), .B1(n17266), .B2(n12554), .ZN(
        n6439) );
  OAI22_X1 U15113 ( .A1(n17273), .A2(n17489), .B1(n17267), .B2(n12553), .ZN(
        n6440) );
  OAI22_X1 U15114 ( .A1(n17273), .A2(n17491), .B1(n17265), .B2(n12552), .ZN(
        n6441) );
  OAI22_X1 U15115 ( .A1(n17274), .A2(n17493), .B1(n17266), .B2(n12551), .ZN(
        n6442) );
  OAI22_X1 U15116 ( .A1(n17274), .A2(n17495), .B1(n17267), .B2(n12550), .ZN(
        n6443) );
  OAI22_X1 U15117 ( .A1(n17274), .A2(n17497), .B1(n17265), .B2(n12549), .ZN(
        n6444) );
  OAI22_X1 U15118 ( .A1(n17274), .A2(n17499), .B1(n17266), .B2(n12548), .ZN(
        n6445) );
  OAI22_X1 U15119 ( .A1(n17274), .A2(n17501), .B1(n17267), .B2(n12547), .ZN(
        n6446) );
  OAI22_X1 U15120 ( .A1(n17275), .A2(n17503), .B1(n17265), .B2(n12546), .ZN(
        n6447) );
  OAI22_X1 U15121 ( .A1(n17275), .A2(n17505), .B1(n13655), .B2(n12545), .ZN(
        n6448) );
  OAI22_X1 U15122 ( .A1(n17275), .A2(n17507), .B1(n17265), .B2(n12544), .ZN(
        n6449) );
  OAI22_X1 U15123 ( .A1(n17275), .A2(n17509), .B1(n13655), .B2(n12543), .ZN(
        n6450) );
  OAI22_X1 U15124 ( .A1(n17275), .A2(n17511), .B1(n17265), .B2(n12542), .ZN(
        n6451) );
  OAI22_X1 U15125 ( .A1(n17276), .A2(n17513), .B1(n13655), .B2(n12541), .ZN(
        n6452) );
  OAI22_X1 U15126 ( .A1(n17276), .A2(n17515), .B1(n17265), .B2(n12540), .ZN(
        n6453) );
  OAI22_X1 U15127 ( .A1(n17276), .A2(n17517), .B1(n17266), .B2(n12539), .ZN(
        n6454) );
  OAI22_X1 U15128 ( .A1(n17276), .A2(n17519), .B1(n17267), .B2(n12538), .ZN(
        n6455) );
  OAI22_X1 U15129 ( .A1(n17276), .A2(n17521), .B1(n17265), .B2(n12537), .ZN(
        n6456) );
  OAI22_X1 U15130 ( .A1(n17277), .A2(n17523), .B1(n17265), .B2(n12536), .ZN(
        n6457) );
  OAI22_X1 U15131 ( .A1(n17277), .A2(n17525), .B1(n17266), .B2(n12535), .ZN(
        n6458) );
  OAI22_X1 U15132 ( .A1(n17277), .A2(n17527), .B1(n17267), .B2(n12534), .ZN(
        n6459) );
  OAI22_X1 U15133 ( .A1(n17277), .A2(n17529), .B1(n17265), .B2(n12533), .ZN(
        n6460) );
  OAI22_X1 U15134 ( .A1(n17277), .A2(n17531), .B1(n17265), .B2(n12532), .ZN(
        n6461) );
  OAI22_X1 U15135 ( .A1(n17278), .A2(n17533), .B1(n13655), .B2(n12531), .ZN(
        n6462) );
  OAI22_X1 U15136 ( .A1(n17278), .A2(n17535), .B1(n17265), .B2(n12530), .ZN(
        n6463) );
  OAI22_X1 U15137 ( .A1(n17278), .A2(n17537), .B1(n13655), .B2(n12529), .ZN(
        n6464) );
  OAI22_X1 U15138 ( .A1(n17278), .A2(n17539), .B1(n17265), .B2(n12528), .ZN(
        n6465) );
  OAI22_X1 U15139 ( .A1(n17278), .A2(n17541), .B1(n13655), .B2(n12527), .ZN(
        n6466) );
  OAI22_X1 U15140 ( .A1(n17279), .A2(n17543), .B1(n17265), .B2(n12526), .ZN(
        n6467) );
  OAI22_X1 U15141 ( .A1(n17279), .A2(n17545), .B1(n13655), .B2(n12525), .ZN(
        n6468) );
  OAI22_X1 U15142 ( .A1(n17279), .A2(n17547), .B1(n17265), .B2(n12524), .ZN(
        n6469) );
  OAI22_X1 U15143 ( .A1(n17279), .A2(n17549), .B1(n13655), .B2(n12523), .ZN(
        n6470) );
  OAI22_X1 U15144 ( .A1(n17279), .A2(n17551), .B1(n17265), .B2(n12522), .ZN(
        n6471) );
  OAI22_X1 U15145 ( .A1(n17289), .A2(n17481), .B1(n17283), .B2(n12493), .ZN(
        n6500) );
  OAI22_X1 U15146 ( .A1(n17290), .A2(n17483), .B1(n17284), .B2(n12492), .ZN(
        n6501) );
  OAI22_X1 U15147 ( .A1(n17290), .A2(n17485), .B1(n17282), .B2(n12491), .ZN(
        n6502) );
  OAI22_X1 U15148 ( .A1(n17290), .A2(n17487), .B1(n17283), .B2(n12490), .ZN(
        n6503) );
  OAI22_X1 U15149 ( .A1(n17290), .A2(n17489), .B1(n17284), .B2(n12489), .ZN(
        n6504) );
  OAI22_X1 U15150 ( .A1(n17290), .A2(n17491), .B1(n17282), .B2(n12488), .ZN(
        n6505) );
  OAI22_X1 U15151 ( .A1(n17291), .A2(n17493), .B1(n17283), .B2(n12487), .ZN(
        n6506) );
  OAI22_X1 U15152 ( .A1(n17291), .A2(n17495), .B1(n17284), .B2(n12486), .ZN(
        n6507) );
  OAI22_X1 U15153 ( .A1(n17291), .A2(n17497), .B1(n17282), .B2(n12485), .ZN(
        n6508) );
  OAI22_X1 U15154 ( .A1(n17291), .A2(n17499), .B1(n17283), .B2(n12484), .ZN(
        n6509) );
  OAI22_X1 U15155 ( .A1(n17291), .A2(n17501), .B1(n17284), .B2(n12483), .ZN(
        n6510) );
  OAI22_X1 U15156 ( .A1(n17292), .A2(n17503), .B1(n17282), .B2(n12482), .ZN(
        n6511) );
  OAI22_X1 U15157 ( .A1(n17292), .A2(n17505), .B1(n13653), .B2(n12481), .ZN(
        n6512) );
  OAI22_X1 U15158 ( .A1(n17292), .A2(n17507), .B1(n17282), .B2(n12480), .ZN(
        n6513) );
  OAI22_X1 U15159 ( .A1(n17292), .A2(n17509), .B1(n13653), .B2(n12479), .ZN(
        n6514) );
  OAI22_X1 U15160 ( .A1(n17292), .A2(n17511), .B1(n17282), .B2(n12478), .ZN(
        n6515) );
  OAI22_X1 U15161 ( .A1(n17293), .A2(n17513), .B1(n13653), .B2(n12477), .ZN(
        n6516) );
  OAI22_X1 U15162 ( .A1(n17293), .A2(n17515), .B1(n17282), .B2(n12476), .ZN(
        n6517) );
  OAI22_X1 U15163 ( .A1(n17293), .A2(n17517), .B1(n17283), .B2(n12475), .ZN(
        n6518) );
  OAI22_X1 U15164 ( .A1(n17293), .A2(n17519), .B1(n17284), .B2(n12474), .ZN(
        n6519) );
  OAI22_X1 U15165 ( .A1(n17293), .A2(n17521), .B1(n17282), .B2(n12473), .ZN(
        n6520) );
  OAI22_X1 U15166 ( .A1(n17294), .A2(n17523), .B1(n17282), .B2(n12472), .ZN(
        n6521) );
  OAI22_X1 U15167 ( .A1(n17294), .A2(n17525), .B1(n17283), .B2(n12471), .ZN(
        n6522) );
  OAI22_X1 U15168 ( .A1(n17294), .A2(n17527), .B1(n17284), .B2(n12470), .ZN(
        n6523) );
  OAI22_X1 U15169 ( .A1(n17294), .A2(n17529), .B1(n17282), .B2(n12469), .ZN(
        n6524) );
  OAI22_X1 U15170 ( .A1(n17294), .A2(n17531), .B1(n17282), .B2(n12468), .ZN(
        n6525) );
  OAI22_X1 U15171 ( .A1(n17295), .A2(n17533), .B1(n13653), .B2(n12467), .ZN(
        n6526) );
  OAI22_X1 U15172 ( .A1(n17295), .A2(n17535), .B1(n17282), .B2(n12466), .ZN(
        n6527) );
  OAI22_X1 U15173 ( .A1(n17295), .A2(n17537), .B1(n13653), .B2(n12465), .ZN(
        n6528) );
  OAI22_X1 U15174 ( .A1(n17295), .A2(n17539), .B1(n17282), .B2(n12464), .ZN(
        n6529) );
  OAI22_X1 U15175 ( .A1(n17295), .A2(n17541), .B1(n13653), .B2(n12463), .ZN(
        n6530) );
  OAI22_X1 U15176 ( .A1(n17296), .A2(n17543), .B1(n17282), .B2(n12462), .ZN(
        n6531) );
  OAI22_X1 U15177 ( .A1(n17296), .A2(n17545), .B1(n13653), .B2(n12461), .ZN(
        n6532) );
  OAI22_X1 U15178 ( .A1(n17296), .A2(n17547), .B1(n17282), .B2(n12460), .ZN(
        n6533) );
  OAI22_X1 U15179 ( .A1(n17296), .A2(n17549), .B1(n13653), .B2(n12459), .ZN(
        n6534) );
  OAI22_X1 U15180 ( .A1(n17296), .A2(n17551), .B1(n17282), .B2(n12458), .ZN(
        n6535) );
  OAI22_X1 U15181 ( .A1(n17097), .A2(n17433), .B1(n7864), .B2(n17095), .ZN(
        n5772) );
  OAI22_X1 U15182 ( .A1(n17097), .A2(n17435), .B1(n7862), .B2(n17095), .ZN(
        n5773) );
  OAI22_X1 U15183 ( .A1(n17097), .A2(n17437), .B1(n7860), .B2(n17095), .ZN(
        n5774) );
  OAI22_X1 U15184 ( .A1(n17097), .A2(n17439), .B1(n7858), .B2(n17095), .ZN(
        n5775) );
  OAI22_X1 U15185 ( .A1(n17097), .A2(n17441), .B1(n7856), .B2(n17095), .ZN(
        n5776) );
  OAI22_X1 U15186 ( .A1(n17098), .A2(n17443), .B1(n7854), .B2(n17095), .ZN(
        n5777) );
  OAI22_X1 U15187 ( .A1(n17098), .A2(n17445), .B1(n7852), .B2(n17095), .ZN(
        n5778) );
  OAI22_X1 U15188 ( .A1(n17098), .A2(n17447), .B1(n7850), .B2(n17095), .ZN(
        n5779) );
  OAI22_X1 U15189 ( .A1(n17098), .A2(n17449), .B1(n7848), .B2(n17095), .ZN(
        n5780) );
  OAI22_X1 U15190 ( .A1(n17098), .A2(n17451), .B1(n7846), .B2(n17095), .ZN(
        n5781) );
  OAI22_X1 U15191 ( .A1(n17099), .A2(n17453), .B1(n7844), .B2(n17095), .ZN(
        n5782) );
  OAI22_X1 U15192 ( .A1(n17099), .A2(n17455), .B1(n7842), .B2(n17095), .ZN(
        n5783) );
  OAI22_X1 U15193 ( .A1(n17099), .A2(n17457), .B1(n7840), .B2(n17096), .ZN(
        n5784) );
  OAI22_X1 U15194 ( .A1(n17099), .A2(n17459), .B1(n7838), .B2(n17096), .ZN(
        n5785) );
  OAI22_X1 U15195 ( .A1(n17099), .A2(n17461), .B1(n7836), .B2(n17096), .ZN(
        n5786) );
  OAI22_X1 U15196 ( .A1(n17100), .A2(n17463), .B1(n7834), .B2(n17096), .ZN(
        n5787) );
  OAI22_X1 U15197 ( .A1(n17100), .A2(n17465), .B1(n7832), .B2(n17096), .ZN(
        n5788) );
  OAI22_X1 U15198 ( .A1(n17100), .A2(n17467), .B1(n7830), .B2(n17096), .ZN(
        n5789) );
  OAI22_X1 U15199 ( .A1(n17100), .A2(n17469), .B1(n7828), .B2(n17096), .ZN(
        n5790) );
  OAI22_X1 U15200 ( .A1(n17100), .A2(n17471), .B1(n7826), .B2(n17096), .ZN(
        n5791) );
  OAI22_X1 U15201 ( .A1(n17101), .A2(n17473), .B1(n7824), .B2(n17096), .ZN(
        n5792) );
  OAI22_X1 U15202 ( .A1(n17101), .A2(n17475), .B1(n7822), .B2(n17096), .ZN(
        n5793) );
  OAI22_X1 U15203 ( .A1(n17101), .A2(n17477), .B1(n7820), .B2(n17096), .ZN(
        n5794) );
  OAI22_X1 U15204 ( .A1(n17101), .A2(n17479), .B1(n7818), .B2(n17096), .ZN(
        n5795) );
  OAI22_X1 U15205 ( .A1(n17101), .A2(n17481), .B1(n7816), .B2(n17095), .ZN(
        n5796) );
  OAI22_X1 U15206 ( .A1(n17102), .A2(n17483), .B1(n7814), .B2(n17096), .ZN(
        n5797) );
  OAI22_X1 U15207 ( .A1(n17102), .A2(n17485), .B1(n7812), .B2(n17094), .ZN(
        n5798) );
  OAI22_X1 U15208 ( .A1(n17102), .A2(n17487), .B1(n7810), .B2(n17095), .ZN(
        n5799) );
  OAI22_X1 U15209 ( .A1(n17102), .A2(n17489), .B1(n7808), .B2(n17096), .ZN(
        n5800) );
  OAI22_X1 U15210 ( .A1(n17102), .A2(n17491), .B1(n7806), .B2(n17094), .ZN(
        n5801) );
  OAI22_X1 U15211 ( .A1(n17103), .A2(n17493), .B1(n7804), .B2(n17095), .ZN(
        n5802) );
  OAI22_X1 U15212 ( .A1(n17103), .A2(n17495), .B1(n7802), .B2(n17096), .ZN(
        n5803) );
  OAI22_X1 U15213 ( .A1(n17103), .A2(n17497), .B1(n7800), .B2(n17094), .ZN(
        n5804) );
  OAI22_X1 U15214 ( .A1(n17103), .A2(n17499), .B1(n7798), .B2(n17095), .ZN(
        n5805) );
  OAI22_X1 U15215 ( .A1(n17103), .A2(n17501), .B1(n7796), .B2(n17096), .ZN(
        n5806) );
  OAI22_X1 U15216 ( .A1(n17104), .A2(n17503), .B1(n7794), .B2(n17094), .ZN(
        n5807) );
  OAI22_X1 U15217 ( .A1(n17104), .A2(n17505), .B1(n7792), .B2(n13666), .ZN(
        n5808) );
  OAI22_X1 U15218 ( .A1(n17104), .A2(n17507), .B1(n7790), .B2(n17094), .ZN(
        n5809) );
  OAI22_X1 U15219 ( .A1(n17104), .A2(n17509), .B1(n7788), .B2(n13666), .ZN(
        n5810) );
  OAI22_X1 U15220 ( .A1(n17104), .A2(n17511), .B1(n7786), .B2(n17094), .ZN(
        n5811) );
  OAI22_X1 U15221 ( .A1(n17105), .A2(n17513), .B1(n7784), .B2(n13666), .ZN(
        n5812) );
  OAI22_X1 U15222 ( .A1(n17105), .A2(n17515), .B1(n7782), .B2(n17094), .ZN(
        n5813) );
  OAI22_X1 U15223 ( .A1(n17105), .A2(n17517), .B1(n7780), .B2(n17095), .ZN(
        n5814) );
  OAI22_X1 U15224 ( .A1(n17105), .A2(n17519), .B1(n7778), .B2(n17096), .ZN(
        n5815) );
  OAI22_X1 U15225 ( .A1(n17105), .A2(n17521), .B1(n7776), .B2(n17094), .ZN(
        n5816) );
  OAI22_X1 U15226 ( .A1(n17106), .A2(n17523), .B1(n7774), .B2(n17094), .ZN(
        n5817) );
  OAI22_X1 U15227 ( .A1(n17106), .A2(n17525), .B1(n7772), .B2(n17095), .ZN(
        n5818) );
  OAI22_X1 U15228 ( .A1(n17106), .A2(n17527), .B1(n7770), .B2(n17096), .ZN(
        n5819) );
  OAI22_X1 U15229 ( .A1(n17106), .A2(n17529), .B1(n7768), .B2(n17094), .ZN(
        n5820) );
  OAI22_X1 U15230 ( .A1(n17106), .A2(n17531), .B1(n7766), .B2(n17094), .ZN(
        n5821) );
  OAI22_X1 U15231 ( .A1(n17107), .A2(n17533), .B1(n7764), .B2(n13666), .ZN(
        n5822) );
  OAI22_X1 U15232 ( .A1(n17107), .A2(n17535), .B1(n7762), .B2(n17094), .ZN(
        n5823) );
  OAI22_X1 U15233 ( .A1(n17107), .A2(n17537), .B1(n7760), .B2(n13666), .ZN(
        n5824) );
  OAI22_X1 U15234 ( .A1(n17107), .A2(n17539), .B1(n7758), .B2(n17094), .ZN(
        n5825) );
  OAI22_X1 U15235 ( .A1(n17107), .A2(n17541), .B1(n7756), .B2(n13666), .ZN(
        n5826) );
  OAI22_X1 U15236 ( .A1(n17108), .A2(n17543), .B1(n7754), .B2(n17094), .ZN(
        n5827) );
  OAI22_X1 U15237 ( .A1(n17108), .A2(n17545), .B1(n7752), .B2(n13666), .ZN(
        n5828) );
  OAI22_X1 U15238 ( .A1(n17108), .A2(n17547), .B1(n7750), .B2(n17094), .ZN(
        n5829) );
  OAI22_X1 U15239 ( .A1(n17108), .A2(n17549), .B1(n7748), .B2(n13666), .ZN(
        n5830) );
  OAI22_X1 U15240 ( .A1(n17108), .A2(n17551), .B1(n7746), .B2(n17094), .ZN(
        n5831) );
  OAI22_X1 U15241 ( .A1(n17109), .A2(n17553), .B1(n7744), .B2(n13666), .ZN(
        n5832) );
  OAI22_X1 U15242 ( .A1(n17109), .A2(n17555), .B1(n7742), .B2(n13666), .ZN(
        n5833) );
  OAI22_X1 U15243 ( .A1(n17109), .A2(n17557), .B1(n7740), .B2(n17094), .ZN(
        n5834) );
  OAI22_X1 U15244 ( .A1(n17109), .A2(n17578), .B1(n7738), .B2(n13666), .ZN(
        n5835) );
  OAI22_X1 U15245 ( .A1(n17114), .A2(n17433), .B1(n7736), .B2(n17112), .ZN(
        n5836) );
  OAI22_X1 U15246 ( .A1(n17114), .A2(n17435), .B1(n7734), .B2(n17112), .ZN(
        n5837) );
  OAI22_X1 U15247 ( .A1(n17114), .A2(n17437), .B1(n7732), .B2(n17112), .ZN(
        n5838) );
  OAI22_X1 U15248 ( .A1(n17114), .A2(n17439), .B1(n7730), .B2(n17112), .ZN(
        n5839) );
  OAI22_X1 U15249 ( .A1(n17114), .A2(n17441), .B1(n7728), .B2(n17112), .ZN(
        n5840) );
  OAI22_X1 U15250 ( .A1(n17115), .A2(n17443), .B1(n7726), .B2(n17112), .ZN(
        n5841) );
  OAI22_X1 U15251 ( .A1(n17115), .A2(n17445), .B1(n7724), .B2(n17112), .ZN(
        n5842) );
  OAI22_X1 U15252 ( .A1(n17115), .A2(n17447), .B1(n7722), .B2(n17112), .ZN(
        n5843) );
  OAI22_X1 U15253 ( .A1(n17115), .A2(n17449), .B1(n7720), .B2(n17112), .ZN(
        n5844) );
  OAI22_X1 U15254 ( .A1(n17115), .A2(n17451), .B1(n7718), .B2(n17112), .ZN(
        n5845) );
  OAI22_X1 U15255 ( .A1(n17116), .A2(n17453), .B1(n7716), .B2(n17112), .ZN(
        n5846) );
  OAI22_X1 U15256 ( .A1(n17116), .A2(n17455), .B1(n7714), .B2(n17112), .ZN(
        n5847) );
  OAI22_X1 U15257 ( .A1(n17116), .A2(n17457), .B1(n7712), .B2(n17113), .ZN(
        n5848) );
  OAI22_X1 U15258 ( .A1(n17116), .A2(n17459), .B1(n7710), .B2(n17113), .ZN(
        n5849) );
  OAI22_X1 U15259 ( .A1(n17116), .A2(n17461), .B1(n7708), .B2(n17113), .ZN(
        n5850) );
  OAI22_X1 U15260 ( .A1(n17117), .A2(n17463), .B1(n7706), .B2(n17113), .ZN(
        n5851) );
  OAI22_X1 U15261 ( .A1(n17117), .A2(n17465), .B1(n7704), .B2(n17113), .ZN(
        n5852) );
  OAI22_X1 U15262 ( .A1(n17117), .A2(n17467), .B1(n7702), .B2(n17113), .ZN(
        n5853) );
  OAI22_X1 U15263 ( .A1(n17117), .A2(n17469), .B1(n7700), .B2(n17113), .ZN(
        n5854) );
  OAI22_X1 U15264 ( .A1(n17117), .A2(n17471), .B1(n7698), .B2(n17113), .ZN(
        n5855) );
  OAI22_X1 U15265 ( .A1(n17118), .A2(n17473), .B1(n7696), .B2(n17113), .ZN(
        n5856) );
  OAI22_X1 U15266 ( .A1(n17118), .A2(n17475), .B1(n7694), .B2(n17113), .ZN(
        n5857) );
  OAI22_X1 U15267 ( .A1(n17118), .A2(n17477), .B1(n7692), .B2(n17113), .ZN(
        n5858) );
  OAI22_X1 U15268 ( .A1(n17118), .A2(n17479), .B1(n7690), .B2(n17113), .ZN(
        n5859) );
  OAI22_X1 U15269 ( .A1(n17118), .A2(n17481), .B1(n7688), .B2(n17112), .ZN(
        n5860) );
  OAI22_X1 U15270 ( .A1(n17119), .A2(n17483), .B1(n7686), .B2(n17113), .ZN(
        n5861) );
  OAI22_X1 U15271 ( .A1(n17119), .A2(n17485), .B1(n7684), .B2(n17111), .ZN(
        n5862) );
  OAI22_X1 U15272 ( .A1(n17119), .A2(n17487), .B1(n7682), .B2(n17112), .ZN(
        n5863) );
  OAI22_X1 U15273 ( .A1(n17119), .A2(n17489), .B1(n7680), .B2(n17113), .ZN(
        n5864) );
  OAI22_X1 U15274 ( .A1(n17119), .A2(n17491), .B1(n7678), .B2(n17111), .ZN(
        n5865) );
  OAI22_X1 U15275 ( .A1(n17120), .A2(n17493), .B1(n7676), .B2(n17112), .ZN(
        n5866) );
  OAI22_X1 U15276 ( .A1(n17120), .A2(n17495), .B1(n7674), .B2(n17113), .ZN(
        n5867) );
  OAI22_X1 U15277 ( .A1(n17120), .A2(n17497), .B1(n7672), .B2(n17111), .ZN(
        n5868) );
  OAI22_X1 U15278 ( .A1(n17120), .A2(n17499), .B1(n7670), .B2(n17112), .ZN(
        n5869) );
  OAI22_X1 U15279 ( .A1(n17120), .A2(n17501), .B1(n7668), .B2(n17113), .ZN(
        n5870) );
  OAI22_X1 U15280 ( .A1(n17121), .A2(n17503), .B1(n7666), .B2(n17111), .ZN(
        n5871) );
  OAI22_X1 U15281 ( .A1(n17121), .A2(n17505), .B1(n7664), .B2(n13665), .ZN(
        n5872) );
  OAI22_X1 U15282 ( .A1(n17121), .A2(n17507), .B1(n7662), .B2(n17111), .ZN(
        n5873) );
  OAI22_X1 U15283 ( .A1(n17121), .A2(n17509), .B1(n7660), .B2(n13665), .ZN(
        n5874) );
  OAI22_X1 U15284 ( .A1(n17121), .A2(n17511), .B1(n7658), .B2(n17111), .ZN(
        n5875) );
  OAI22_X1 U15285 ( .A1(n17122), .A2(n17513), .B1(n7656), .B2(n13665), .ZN(
        n5876) );
  OAI22_X1 U15286 ( .A1(n17122), .A2(n17515), .B1(n7654), .B2(n17111), .ZN(
        n5877) );
  OAI22_X1 U15287 ( .A1(n17122), .A2(n17517), .B1(n7652), .B2(n17112), .ZN(
        n5878) );
  OAI22_X1 U15288 ( .A1(n17122), .A2(n17519), .B1(n7650), .B2(n17113), .ZN(
        n5879) );
  OAI22_X1 U15289 ( .A1(n17122), .A2(n17521), .B1(n7648), .B2(n17111), .ZN(
        n5880) );
  OAI22_X1 U15290 ( .A1(n17123), .A2(n17523), .B1(n7646), .B2(n17111), .ZN(
        n5881) );
  OAI22_X1 U15291 ( .A1(n17123), .A2(n17525), .B1(n7644), .B2(n17112), .ZN(
        n5882) );
  OAI22_X1 U15292 ( .A1(n17123), .A2(n17527), .B1(n7642), .B2(n17113), .ZN(
        n5883) );
  OAI22_X1 U15293 ( .A1(n17123), .A2(n17529), .B1(n7640), .B2(n17111), .ZN(
        n5884) );
  OAI22_X1 U15294 ( .A1(n17123), .A2(n17531), .B1(n7638), .B2(n17111), .ZN(
        n5885) );
  OAI22_X1 U15295 ( .A1(n17124), .A2(n17533), .B1(n7636), .B2(n13665), .ZN(
        n5886) );
  OAI22_X1 U15296 ( .A1(n17124), .A2(n17535), .B1(n7634), .B2(n17111), .ZN(
        n5887) );
  OAI22_X1 U15297 ( .A1(n17124), .A2(n17537), .B1(n7632), .B2(n13665), .ZN(
        n5888) );
  OAI22_X1 U15298 ( .A1(n17124), .A2(n17539), .B1(n7630), .B2(n17111), .ZN(
        n5889) );
  OAI22_X1 U15299 ( .A1(n17124), .A2(n17541), .B1(n7628), .B2(n13665), .ZN(
        n5890) );
  OAI22_X1 U15300 ( .A1(n17125), .A2(n17543), .B1(n7626), .B2(n17111), .ZN(
        n5891) );
  OAI22_X1 U15301 ( .A1(n17125), .A2(n17545), .B1(n7624), .B2(n13665), .ZN(
        n5892) );
  OAI22_X1 U15302 ( .A1(n17125), .A2(n17547), .B1(n7622), .B2(n17111), .ZN(
        n5893) );
  OAI22_X1 U15303 ( .A1(n17125), .A2(n17549), .B1(n7620), .B2(n13665), .ZN(
        n5894) );
  OAI22_X1 U15304 ( .A1(n17125), .A2(n17551), .B1(n7618), .B2(n17111), .ZN(
        n5895) );
  OAI22_X1 U15305 ( .A1(n17126), .A2(n17553), .B1(n7616), .B2(n13665), .ZN(
        n5896) );
  OAI22_X1 U15306 ( .A1(n17126), .A2(n17555), .B1(n7614), .B2(n13665), .ZN(
        n5897) );
  OAI22_X1 U15307 ( .A1(n17126), .A2(n17557), .B1(n7612), .B2(n17111), .ZN(
        n5898) );
  OAI22_X1 U15308 ( .A1(n17126), .A2(n17578), .B1(n7610), .B2(n13665), .ZN(
        n5899) );
  OAI22_X1 U15309 ( .A1(n17200), .A2(n17433), .B1(n900), .B2(n17198), .ZN(
        n6156) );
  OAI22_X1 U15310 ( .A1(n17200), .A2(n17435), .B1(n899), .B2(n17198), .ZN(
        n6157) );
  OAI22_X1 U15311 ( .A1(n17200), .A2(n17437), .B1(n898), .B2(n17198), .ZN(
        n6158) );
  OAI22_X1 U15312 ( .A1(n17200), .A2(n17439), .B1(n897), .B2(n17198), .ZN(
        n6159) );
  OAI22_X1 U15313 ( .A1(n17200), .A2(n17441), .B1(n896), .B2(n17198), .ZN(
        n6160) );
  OAI22_X1 U15314 ( .A1(n17201), .A2(n17443), .B1(n895), .B2(n17198), .ZN(
        n6161) );
  OAI22_X1 U15315 ( .A1(n17201), .A2(n17445), .B1(n894), .B2(n17198), .ZN(
        n6162) );
  OAI22_X1 U15316 ( .A1(n17201), .A2(n17447), .B1(n893), .B2(n17198), .ZN(
        n6163) );
  OAI22_X1 U15317 ( .A1(n17201), .A2(n17449), .B1(n892), .B2(n17198), .ZN(
        n6164) );
  OAI22_X1 U15318 ( .A1(n17201), .A2(n17451), .B1(n891), .B2(n17198), .ZN(
        n6165) );
  OAI22_X1 U15319 ( .A1(n17202), .A2(n17453), .B1(n890), .B2(n17198), .ZN(
        n6166) );
  OAI22_X1 U15320 ( .A1(n17202), .A2(n17455), .B1(n889), .B2(n17198), .ZN(
        n6167) );
  OAI22_X1 U15321 ( .A1(n17202), .A2(n17457), .B1(n888), .B2(n17199), .ZN(
        n6168) );
  OAI22_X1 U15322 ( .A1(n17202), .A2(n17459), .B1(n887), .B2(n17199), .ZN(
        n6169) );
  OAI22_X1 U15323 ( .A1(n17202), .A2(n17461), .B1(n886), .B2(n17199), .ZN(
        n6170) );
  OAI22_X1 U15324 ( .A1(n17203), .A2(n17463), .B1(n885), .B2(n17199), .ZN(
        n6171) );
  OAI22_X1 U15325 ( .A1(n17203), .A2(n17465), .B1(n884), .B2(n17199), .ZN(
        n6172) );
  OAI22_X1 U15326 ( .A1(n17203), .A2(n17467), .B1(n883), .B2(n17199), .ZN(
        n6173) );
  OAI22_X1 U15327 ( .A1(n17203), .A2(n17469), .B1(n882), .B2(n17199), .ZN(
        n6174) );
  OAI22_X1 U15328 ( .A1(n17203), .A2(n17471), .B1(n881), .B2(n17199), .ZN(
        n6175) );
  OAI22_X1 U15329 ( .A1(n17204), .A2(n17473), .B1(n880), .B2(n17199), .ZN(
        n6176) );
  OAI22_X1 U15330 ( .A1(n17204), .A2(n17475), .B1(n879), .B2(n17199), .ZN(
        n6177) );
  OAI22_X1 U15331 ( .A1(n17204), .A2(n17477), .B1(n878), .B2(n17199), .ZN(
        n6178) );
  OAI22_X1 U15332 ( .A1(n17204), .A2(n17479), .B1(n877), .B2(n17199), .ZN(
        n6179) );
  OAI22_X1 U15333 ( .A1(n17204), .A2(n17481), .B1(n876), .B2(n17198), .ZN(
        n6180) );
  OAI22_X1 U15334 ( .A1(n17205), .A2(n17483), .B1(n875), .B2(n17199), .ZN(
        n6181) );
  OAI22_X1 U15335 ( .A1(n17205), .A2(n17485), .B1(n874), .B2(n17197), .ZN(
        n6182) );
  OAI22_X1 U15336 ( .A1(n17205), .A2(n17487), .B1(n873), .B2(n17198), .ZN(
        n6183) );
  OAI22_X1 U15337 ( .A1(n17205), .A2(n17489), .B1(n872), .B2(n17199), .ZN(
        n6184) );
  OAI22_X1 U15338 ( .A1(n17205), .A2(n17491), .B1(n871), .B2(n17197), .ZN(
        n6185) );
  OAI22_X1 U15339 ( .A1(n17206), .A2(n17493), .B1(n870), .B2(n17198), .ZN(
        n6186) );
  OAI22_X1 U15340 ( .A1(n17206), .A2(n17495), .B1(n869), .B2(n17199), .ZN(
        n6187) );
  OAI22_X1 U15341 ( .A1(n17206), .A2(n17497), .B1(n868), .B2(n17197), .ZN(
        n6188) );
  OAI22_X1 U15342 ( .A1(n17206), .A2(n17499), .B1(n867), .B2(n17198), .ZN(
        n6189) );
  OAI22_X1 U15343 ( .A1(n17206), .A2(n17501), .B1(n866), .B2(n17199), .ZN(
        n6190) );
  OAI22_X1 U15344 ( .A1(n17207), .A2(n17503), .B1(n865), .B2(n17197), .ZN(
        n6191) );
  OAI22_X1 U15345 ( .A1(n17207), .A2(n17505), .B1(n864), .B2(n13659), .ZN(
        n6192) );
  OAI22_X1 U15346 ( .A1(n17207), .A2(n17507), .B1(n863), .B2(n17197), .ZN(
        n6193) );
  OAI22_X1 U15347 ( .A1(n17207), .A2(n17509), .B1(n862), .B2(n13659), .ZN(
        n6194) );
  OAI22_X1 U15348 ( .A1(n17207), .A2(n17511), .B1(n861), .B2(n17197), .ZN(
        n6195) );
  OAI22_X1 U15349 ( .A1(n17208), .A2(n17513), .B1(n860), .B2(n13659), .ZN(
        n6196) );
  OAI22_X1 U15350 ( .A1(n17208), .A2(n17515), .B1(n859), .B2(n17197), .ZN(
        n6197) );
  OAI22_X1 U15351 ( .A1(n17208), .A2(n17517), .B1(n858), .B2(n17198), .ZN(
        n6198) );
  OAI22_X1 U15352 ( .A1(n17208), .A2(n17519), .B1(n857), .B2(n17199), .ZN(
        n6199) );
  OAI22_X1 U15353 ( .A1(n17208), .A2(n17521), .B1(n856), .B2(n17197), .ZN(
        n6200) );
  OAI22_X1 U15354 ( .A1(n17209), .A2(n17523), .B1(n855), .B2(n17197), .ZN(
        n6201) );
  OAI22_X1 U15355 ( .A1(n17209), .A2(n17525), .B1(n854), .B2(n17198), .ZN(
        n6202) );
  OAI22_X1 U15356 ( .A1(n17209), .A2(n17527), .B1(n853), .B2(n17199), .ZN(
        n6203) );
  OAI22_X1 U15357 ( .A1(n17209), .A2(n17529), .B1(n852), .B2(n17197), .ZN(
        n6204) );
  OAI22_X1 U15358 ( .A1(n17209), .A2(n17531), .B1(n851), .B2(n17197), .ZN(
        n6205) );
  OAI22_X1 U15359 ( .A1(n17210), .A2(n17533), .B1(n850), .B2(n13659), .ZN(
        n6206) );
  OAI22_X1 U15360 ( .A1(n17210), .A2(n17535), .B1(n849), .B2(n17197), .ZN(
        n6207) );
  OAI22_X1 U15361 ( .A1(n17210), .A2(n17537), .B1(n848), .B2(n13659), .ZN(
        n6208) );
  OAI22_X1 U15362 ( .A1(n17210), .A2(n17539), .B1(n847), .B2(n17197), .ZN(
        n6209) );
  OAI22_X1 U15363 ( .A1(n17210), .A2(n17541), .B1(n846), .B2(n13659), .ZN(
        n6210) );
  OAI22_X1 U15364 ( .A1(n17211), .A2(n17543), .B1(n845), .B2(n17197), .ZN(
        n6211) );
  OAI22_X1 U15365 ( .A1(n17211), .A2(n17545), .B1(n844), .B2(n13659), .ZN(
        n6212) );
  OAI22_X1 U15366 ( .A1(n17211), .A2(n17547), .B1(n843), .B2(n17197), .ZN(
        n6213) );
  OAI22_X1 U15367 ( .A1(n17211), .A2(n17549), .B1(n842), .B2(n13659), .ZN(
        n6214) );
  OAI22_X1 U15368 ( .A1(n17211), .A2(n17551), .B1(n841), .B2(n17197), .ZN(
        n6215) );
  OAI22_X1 U15369 ( .A1(n17212), .A2(n17553), .B1(n840), .B2(n13659), .ZN(
        n6216) );
  OAI22_X1 U15370 ( .A1(n17212), .A2(n17555), .B1(n839), .B2(n13659), .ZN(
        n6217) );
  OAI22_X1 U15371 ( .A1(n17212), .A2(n17557), .B1(n838), .B2(n17197), .ZN(
        n6218) );
  OAI22_X1 U15372 ( .A1(n17212), .A2(n17578), .B1(n837), .B2(n13659), .ZN(
        n6219) );
  OAI22_X1 U15373 ( .A1(n17303), .A2(n17432), .B1(n16413), .B2(n17300), .ZN(
        n6540) );
  OAI22_X1 U15374 ( .A1(n17303), .A2(n17434), .B1(n16408), .B2(n17300), .ZN(
        n6541) );
  OAI22_X1 U15375 ( .A1(n17303), .A2(n17436), .B1(n16403), .B2(n17300), .ZN(
        n6542) );
  OAI22_X1 U15376 ( .A1(n17303), .A2(n17438), .B1(n16398), .B2(n17300), .ZN(
        n6543) );
  OAI22_X1 U15377 ( .A1(n17303), .A2(n17440), .B1(n16393), .B2(n17300), .ZN(
        n6544) );
  OAI22_X1 U15378 ( .A1(n17304), .A2(n17442), .B1(n16388), .B2(n17300), .ZN(
        n6545) );
  OAI22_X1 U15379 ( .A1(n17304), .A2(n17444), .B1(n16383), .B2(n17300), .ZN(
        n6546) );
  OAI22_X1 U15380 ( .A1(n17304), .A2(n17446), .B1(n16378), .B2(n17300), .ZN(
        n6547) );
  OAI22_X1 U15381 ( .A1(n17304), .A2(n17448), .B1(n16373), .B2(n17300), .ZN(
        n6548) );
  OAI22_X1 U15382 ( .A1(n17304), .A2(n17450), .B1(n16368), .B2(n17300), .ZN(
        n6549) );
  OAI22_X1 U15383 ( .A1(n17305), .A2(n17452), .B1(n16363), .B2(n17300), .ZN(
        n6550) );
  OAI22_X1 U15384 ( .A1(n17305), .A2(n17454), .B1(n16358), .B2(n17300), .ZN(
        n6551) );
  OAI22_X1 U15385 ( .A1(n17305), .A2(n17456), .B1(n16353), .B2(n17301), .ZN(
        n6552) );
  OAI22_X1 U15386 ( .A1(n17305), .A2(n17458), .B1(n16348), .B2(n17301), .ZN(
        n6553) );
  OAI22_X1 U15387 ( .A1(n17305), .A2(n17460), .B1(n16343), .B2(n17301), .ZN(
        n6554) );
  OAI22_X1 U15388 ( .A1(n17306), .A2(n17462), .B1(n16338), .B2(n17301), .ZN(
        n6555) );
  OAI22_X1 U15389 ( .A1(n17306), .A2(n17464), .B1(n16333), .B2(n17301), .ZN(
        n6556) );
  OAI22_X1 U15390 ( .A1(n17306), .A2(n17466), .B1(n16328), .B2(n17301), .ZN(
        n6557) );
  OAI22_X1 U15391 ( .A1(n17306), .A2(n17468), .B1(n16323), .B2(n17301), .ZN(
        n6558) );
  OAI22_X1 U15392 ( .A1(n17306), .A2(n17470), .B1(n16318), .B2(n17301), .ZN(
        n6559) );
  OAI22_X1 U15393 ( .A1(n17307), .A2(n17472), .B1(n16313), .B2(n17301), .ZN(
        n6560) );
  OAI22_X1 U15394 ( .A1(n17307), .A2(n17474), .B1(n16308), .B2(n17301), .ZN(
        n6561) );
  OAI22_X1 U15395 ( .A1(n17307), .A2(n17476), .B1(n16303), .B2(n17301), .ZN(
        n6562) );
  OAI22_X1 U15396 ( .A1(n17307), .A2(n17478), .B1(n16298), .B2(n17301), .ZN(
        n6563) );
  OAI22_X1 U15397 ( .A1(n17307), .A2(n17480), .B1(n16293), .B2(n17302), .ZN(
        n6564) );
  OAI22_X1 U15398 ( .A1(n17308), .A2(n17482), .B1(n16288), .B2(n17302), .ZN(
        n6565) );
  OAI22_X1 U15399 ( .A1(n17308), .A2(n17484), .B1(n16283), .B2(n17302), .ZN(
        n6566) );
  OAI22_X1 U15400 ( .A1(n17308), .A2(n17486), .B1(n16278), .B2(n17302), .ZN(
        n6567) );
  OAI22_X1 U15401 ( .A1(n17308), .A2(n17488), .B1(n16273), .B2(n17302), .ZN(
        n6568) );
  OAI22_X1 U15402 ( .A1(n17308), .A2(n17490), .B1(n16268), .B2(n17302), .ZN(
        n6569) );
  OAI22_X1 U15403 ( .A1(n17309), .A2(n17492), .B1(n16263), .B2(n17302), .ZN(
        n6570) );
  OAI22_X1 U15404 ( .A1(n17309), .A2(n17494), .B1(n16258), .B2(n17302), .ZN(
        n6571) );
  OAI22_X1 U15405 ( .A1(n17309), .A2(n17496), .B1(n16253), .B2(n17302), .ZN(
        n6572) );
  OAI22_X1 U15406 ( .A1(n17309), .A2(n17498), .B1(n16248), .B2(n17302), .ZN(
        n6573) );
  OAI22_X1 U15407 ( .A1(n17309), .A2(n17500), .B1(n16243), .B2(n17302), .ZN(
        n6574) );
  OAI22_X1 U15408 ( .A1(n17310), .A2(n17502), .B1(n16238), .B2(n17302), .ZN(
        n6575) );
  OAI22_X1 U15409 ( .A1(n17310), .A2(n17504), .B1(n16233), .B2(n13650), .ZN(
        n6576) );
  OAI22_X1 U15410 ( .A1(n17310), .A2(n17506), .B1(n16228), .B2(n17299), .ZN(
        n6577) );
  OAI22_X1 U15411 ( .A1(n17310), .A2(n17508), .B1(n16223), .B2(n13650), .ZN(
        n6578) );
  OAI22_X1 U15412 ( .A1(n17310), .A2(n17510), .B1(n16218), .B2(n17299), .ZN(
        n6579) );
  OAI22_X1 U15413 ( .A1(n17311), .A2(n17512), .B1(n16213), .B2(n13650), .ZN(
        n6580) );
  OAI22_X1 U15414 ( .A1(n17311), .A2(n17514), .B1(n16208), .B2(n17299), .ZN(
        n6581) );
  OAI22_X1 U15415 ( .A1(n17311), .A2(n17516), .B1(n16203), .B2(n17300), .ZN(
        n6582) );
  OAI22_X1 U15416 ( .A1(n17311), .A2(n17518), .B1(n16198), .B2(n17301), .ZN(
        n6583) );
  OAI22_X1 U15417 ( .A1(n17311), .A2(n17520), .B1(n16193), .B2(n17302), .ZN(
        n6584) );
  OAI22_X1 U15418 ( .A1(n17312), .A2(n17522), .B1(n16188), .B2(n17299), .ZN(
        n6585) );
  OAI22_X1 U15419 ( .A1(n17312), .A2(n17524), .B1(n16183), .B2(n17300), .ZN(
        n6586) );
  OAI22_X1 U15420 ( .A1(n17312), .A2(n17526), .B1(n16178), .B2(n17301), .ZN(
        n6587) );
  OAI22_X1 U15421 ( .A1(n17312), .A2(n17528), .B1(n16173), .B2(n17299), .ZN(
        n6588) );
  OAI22_X1 U15422 ( .A1(n17312), .A2(n17530), .B1(n16168), .B2(n17299), .ZN(
        n6589) );
  OAI22_X1 U15423 ( .A1(n17313), .A2(n17532), .B1(n16163), .B2(n13650), .ZN(
        n6590) );
  OAI22_X1 U15424 ( .A1(n17313), .A2(n17534), .B1(n16158), .B2(n17299), .ZN(
        n6591) );
  OAI22_X1 U15425 ( .A1(n17313), .A2(n17536), .B1(n16153), .B2(n13650), .ZN(
        n6592) );
  OAI22_X1 U15426 ( .A1(n17313), .A2(n17538), .B1(n16148), .B2(n17299), .ZN(
        n6593) );
  OAI22_X1 U15427 ( .A1(n17313), .A2(n17540), .B1(n16143), .B2(n13650), .ZN(
        n6594) );
  OAI22_X1 U15428 ( .A1(n17314), .A2(n17542), .B1(n16138), .B2(n17299), .ZN(
        n6595) );
  OAI22_X1 U15429 ( .A1(n17314), .A2(n17544), .B1(n16133), .B2(n13650), .ZN(
        n6596) );
  OAI22_X1 U15430 ( .A1(n17314), .A2(n17546), .B1(n16128), .B2(n17299), .ZN(
        n6597) );
  OAI22_X1 U15431 ( .A1(n17314), .A2(n17548), .B1(n16123), .B2(n13650), .ZN(
        n6598) );
  OAI22_X1 U15432 ( .A1(n17314), .A2(n17550), .B1(n16118), .B2(n17299), .ZN(
        n6599) );
  OAI22_X1 U15433 ( .A1(n17315), .A2(n17552), .B1(n16113), .B2(n13650), .ZN(
        n6600) );
  OAI22_X1 U15434 ( .A1(n17315), .A2(n17554), .B1(n16108), .B2(n13650), .ZN(
        n6601) );
  OAI22_X1 U15435 ( .A1(n17315), .A2(n17556), .B1(n16103), .B2(n17299), .ZN(
        n6602) );
  OAI22_X1 U15436 ( .A1(n17315), .A2(n17577), .B1(n16098), .B2(n13650), .ZN(
        n6603) );
  OAI22_X1 U15437 ( .A1(n17398), .A2(n17433), .B1(n16411), .B2(n17395), .ZN(
        n6860) );
  OAI22_X1 U15438 ( .A1(n17398), .A2(n17435), .B1(n16406), .B2(n17395), .ZN(
        n6861) );
  OAI22_X1 U15439 ( .A1(n17398), .A2(n17437), .B1(n16401), .B2(n17395), .ZN(
        n6862) );
  OAI22_X1 U15440 ( .A1(n17398), .A2(n17439), .B1(n16396), .B2(n17395), .ZN(
        n6863) );
  OAI22_X1 U15441 ( .A1(n17398), .A2(n17441), .B1(n16391), .B2(n17395), .ZN(
        n6864) );
  OAI22_X1 U15442 ( .A1(n17399), .A2(n17443), .B1(n16386), .B2(n17395), .ZN(
        n6865) );
  OAI22_X1 U15443 ( .A1(n17399), .A2(n17445), .B1(n16381), .B2(n17395), .ZN(
        n6866) );
  OAI22_X1 U15444 ( .A1(n17399), .A2(n17447), .B1(n16376), .B2(n17395), .ZN(
        n6867) );
  OAI22_X1 U15445 ( .A1(n17399), .A2(n17449), .B1(n16371), .B2(n17395), .ZN(
        n6868) );
  OAI22_X1 U15446 ( .A1(n17399), .A2(n17451), .B1(n16366), .B2(n17395), .ZN(
        n6869) );
  OAI22_X1 U15447 ( .A1(n17400), .A2(n17453), .B1(n16361), .B2(n17395), .ZN(
        n6870) );
  OAI22_X1 U15448 ( .A1(n17400), .A2(n17455), .B1(n16356), .B2(n17395), .ZN(
        n6871) );
  OAI22_X1 U15449 ( .A1(n17400), .A2(n17457), .B1(n16351), .B2(n17396), .ZN(
        n6872) );
  OAI22_X1 U15450 ( .A1(n17400), .A2(n17459), .B1(n16346), .B2(n17396), .ZN(
        n6873) );
  OAI22_X1 U15451 ( .A1(n17400), .A2(n17461), .B1(n16341), .B2(n17396), .ZN(
        n6874) );
  OAI22_X1 U15452 ( .A1(n17401), .A2(n17463), .B1(n16336), .B2(n17396), .ZN(
        n6875) );
  OAI22_X1 U15453 ( .A1(n17401), .A2(n17465), .B1(n16331), .B2(n17396), .ZN(
        n6876) );
  OAI22_X1 U15454 ( .A1(n17401), .A2(n17467), .B1(n16326), .B2(n17396), .ZN(
        n6877) );
  OAI22_X1 U15455 ( .A1(n17401), .A2(n17469), .B1(n16321), .B2(n17396), .ZN(
        n6878) );
  OAI22_X1 U15456 ( .A1(n17401), .A2(n17471), .B1(n16316), .B2(n17396), .ZN(
        n6879) );
  OAI22_X1 U15457 ( .A1(n17402), .A2(n17473), .B1(n16311), .B2(n17396), .ZN(
        n6880) );
  OAI22_X1 U15458 ( .A1(n17402), .A2(n17475), .B1(n16306), .B2(n17396), .ZN(
        n6881) );
  OAI22_X1 U15459 ( .A1(n17402), .A2(n17477), .B1(n16301), .B2(n17396), .ZN(
        n6882) );
  OAI22_X1 U15460 ( .A1(n17402), .A2(n17479), .B1(n16296), .B2(n17396), .ZN(
        n6883) );
  OAI22_X1 U15461 ( .A1(n17402), .A2(n17481), .B1(n16291), .B2(n17397), .ZN(
        n6884) );
  OAI22_X1 U15462 ( .A1(n17403), .A2(n17483), .B1(n16286), .B2(n17397), .ZN(
        n6885) );
  OAI22_X1 U15463 ( .A1(n17403), .A2(n17485), .B1(n16281), .B2(n17397), .ZN(
        n6886) );
  OAI22_X1 U15464 ( .A1(n17403), .A2(n17487), .B1(n16276), .B2(n17397), .ZN(
        n6887) );
  OAI22_X1 U15465 ( .A1(n17403), .A2(n17489), .B1(n16271), .B2(n17397), .ZN(
        n6888) );
  OAI22_X1 U15466 ( .A1(n17403), .A2(n17491), .B1(n16266), .B2(n17397), .ZN(
        n6889) );
  OAI22_X1 U15467 ( .A1(n17404), .A2(n17493), .B1(n16261), .B2(n17397), .ZN(
        n6890) );
  OAI22_X1 U15468 ( .A1(n17404), .A2(n17495), .B1(n16256), .B2(n17397), .ZN(
        n6891) );
  OAI22_X1 U15469 ( .A1(n17404), .A2(n17497), .B1(n16251), .B2(n17397), .ZN(
        n6892) );
  OAI22_X1 U15470 ( .A1(n17404), .A2(n17499), .B1(n16246), .B2(n17397), .ZN(
        n6893) );
  OAI22_X1 U15471 ( .A1(n17404), .A2(n17501), .B1(n16241), .B2(n17397), .ZN(
        n6894) );
  OAI22_X1 U15472 ( .A1(n17405), .A2(n17503), .B1(n16236), .B2(n17397), .ZN(
        n6895) );
  OAI22_X1 U15473 ( .A1(n17405), .A2(n17505), .B1(n16231), .B2(n13640), .ZN(
        n6896) );
  OAI22_X1 U15474 ( .A1(n17405), .A2(n17507), .B1(n16226), .B2(n17394), .ZN(
        n6897) );
  OAI22_X1 U15475 ( .A1(n17405), .A2(n17509), .B1(n16221), .B2(n13640), .ZN(
        n6898) );
  OAI22_X1 U15476 ( .A1(n17405), .A2(n17511), .B1(n16216), .B2(n17394), .ZN(
        n6899) );
  OAI22_X1 U15477 ( .A1(n17406), .A2(n17513), .B1(n16211), .B2(n13640), .ZN(
        n6900) );
  OAI22_X1 U15478 ( .A1(n17406), .A2(n17515), .B1(n16206), .B2(n17394), .ZN(
        n6901) );
  OAI22_X1 U15479 ( .A1(n17406), .A2(n17517), .B1(n16201), .B2(n17395), .ZN(
        n6902) );
  OAI22_X1 U15480 ( .A1(n17406), .A2(n17519), .B1(n16196), .B2(n17396), .ZN(
        n6903) );
  OAI22_X1 U15481 ( .A1(n17406), .A2(n17521), .B1(n16191), .B2(n17397), .ZN(
        n6904) );
  OAI22_X1 U15482 ( .A1(n17407), .A2(n17523), .B1(n16186), .B2(n17394), .ZN(
        n6905) );
  OAI22_X1 U15483 ( .A1(n17407), .A2(n17525), .B1(n16181), .B2(n17395), .ZN(
        n6906) );
  OAI22_X1 U15484 ( .A1(n17407), .A2(n17527), .B1(n16176), .B2(n17396), .ZN(
        n6907) );
  OAI22_X1 U15485 ( .A1(n17407), .A2(n17529), .B1(n16171), .B2(n17394), .ZN(
        n6908) );
  OAI22_X1 U15486 ( .A1(n17407), .A2(n17531), .B1(n16166), .B2(n17394), .ZN(
        n6909) );
  OAI22_X1 U15487 ( .A1(n17408), .A2(n17533), .B1(n16161), .B2(n13640), .ZN(
        n6910) );
  OAI22_X1 U15488 ( .A1(n17408), .A2(n17535), .B1(n16156), .B2(n17394), .ZN(
        n6911) );
  OAI22_X1 U15489 ( .A1(n17408), .A2(n17537), .B1(n16151), .B2(n13640), .ZN(
        n6912) );
  OAI22_X1 U15490 ( .A1(n17408), .A2(n17539), .B1(n16146), .B2(n17394), .ZN(
        n6913) );
  OAI22_X1 U15491 ( .A1(n17408), .A2(n17541), .B1(n16141), .B2(n13640), .ZN(
        n6914) );
  OAI22_X1 U15492 ( .A1(n17409), .A2(n17543), .B1(n16136), .B2(n17394), .ZN(
        n6915) );
  OAI22_X1 U15493 ( .A1(n17409), .A2(n17545), .B1(n16131), .B2(n13640), .ZN(
        n6916) );
  OAI22_X1 U15494 ( .A1(n17409), .A2(n17547), .B1(n16126), .B2(n17394), .ZN(
        n6917) );
  OAI22_X1 U15495 ( .A1(n17409), .A2(n17549), .B1(n16121), .B2(n13640), .ZN(
        n6918) );
  OAI22_X1 U15496 ( .A1(n17409), .A2(n17551), .B1(n16116), .B2(n17394), .ZN(
        n6919) );
  OAI22_X1 U15497 ( .A1(n17410), .A2(n17553), .B1(n16111), .B2(n13640), .ZN(
        n6920) );
  OAI22_X1 U15498 ( .A1(n17410), .A2(n17555), .B1(n16106), .B2(n13640), .ZN(
        n6921) );
  OAI22_X1 U15499 ( .A1(n17410), .A2(n17557), .B1(n16101), .B2(n17394), .ZN(
        n6922) );
  OAI22_X1 U15500 ( .A1(n17410), .A2(n17578), .B1(n16096), .B2(n13640), .ZN(
        n6923) );
  OAI22_X1 U15501 ( .A1(n16927), .A2(n17432), .B1(n7863), .B2(n16925), .ZN(
        n5132) );
  OAI22_X1 U15502 ( .A1(n16927), .A2(n17434), .B1(n7861), .B2(n16925), .ZN(
        n5133) );
  OAI22_X1 U15503 ( .A1(n16927), .A2(n17436), .B1(n7859), .B2(n16925), .ZN(
        n5134) );
  OAI22_X1 U15504 ( .A1(n16927), .A2(n17438), .B1(n7857), .B2(n16925), .ZN(
        n5135) );
  OAI22_X1 U15505 ( .A1(n16927), .A2(n17440), .B1(n7855), .B2(n16925), .ZN(
        n5136) );
  OAI22_X1 U15506 ( .A1(n16928), .A2(n17442), .B1(n7853), .B2(n16925), .ZN(
        n5137) );
  OAI22_X1 U15507 ( .A1(n16928), .A2(n17444), .B1(n7851), .B2(n16925), .ZN(
        n5138) );
  OAI22_X1 U15508 ( .A1(n16928), .A2(n17446), .B1(n7849), .B2(n16925), .ZN(
        n5139) );
  OAI22_X1 U15509 ( .A1(n16928), .A2(n17448), .B1(n7847), .B2(n16925), .ZN(
        n5140) );
  OAI22_X1 U15510 ( .A1(n16928), .A2(n17450), .B1(n7845), .B2(n16925), .ZN(
        n5141) );
  OAI22_X1 U15511 ( .A1(n16929), .A2(n17452), .B1(n7843), .B2(n16925), .ZN(
        n5142) );
  OAI22_X1 U15512 ( .A1(n16929), .A2(n17454), .B1(n7841), .B2(n16925), .ZN(
        n5143) );
  OAI22_X1 U15513 ( .A1(n16929), .A2(n17456), .B1(n7839), .B2(n16926), .ZN(
        n5144) );
  OAI22_X1 U15514 ( .A1(n16929), .A2(n17458), .B1(n7837), .B2(n16926), .ZN(
        n5145) );
  OAI22_X1 U15515 ( .A1(n16929), .A2(n17460), .B1(n7835), .B2(n16926), .ZN(
        n5146) );
  OAI22_X1 U15516 ( .A1(n16930), .A2(n17462), .B1(n7833), .B2(n16926), .ZN(
        n5147) );
  OAI22_X1 U15517 ( .A1(n16930), .A2(n17464), .B1(n7831), .B2(n16926), .ZN(
        n5148) );
  OAI22_X1 U15518 ( .A1(n16930), .A2(n17466), .B1(n7829), .B2(n16926), .ZN(
        n5149) );
  OAI22_X1 U15519 ( .A1(n16930), .A2(n17468), .B1(n7827), .B2(n16926), .ZN(
        n5150) );
  OAI22_X1 U15520 ( .A1(n16930), .A2(n17470), .B1(n7825), .B2(n16926), .ZN(
        n5151) );
  OAI22_X1 U15521 ( .A1(n16931), .A2(n17472), .B1(n7823), .B2(n16926), .ZN(
        n5152) );
  OAI22_X1 U15522 ( .A1(n16931), .A2(n17474), .B1(n7821), .B2(n16926), .ZN(
        n5153) );
  OAI22_X1 U15523 ( .A1(n16931), .A2(n17476), .B1(n7819), .B2(n16926), .ZN(
        n5154) );
  OAI22_X1 U15524 ( .A1(n16931), .A2(n17478), .B1(n7817), .B2(n16926), .ZN(
        n5155) );
  OAI22_X1 U15525 ( .A1(n16944), .A2(n17432), .B1(n7735), .B2(n16942), .ZN(
        n5196) );
  OAI22_X1 U15526 ( .A1(n16944), .A2(n17434), .B1(n7733), .B2(n16942), .ZN(
        n5197) );
  OAI22_X1 U15527 ( .A1(n16944), .A2(n17436), .B1(n7731), .B2(n16942), .ZN(
        n5198) );
  OAI22_X1 U15528 ( .A1(n16944), .A2(n17438), .B1(n7729), .B2(n16942), .ZN(
        n5199) );
  OAI22_X1 U15529 ( .A1(n16944), .A2(n17440), .B1(n7727), .B2(n16942), .ZN(
        n5200) );
  OAI22_X1 U15530 ( .A1(n16945), .A2(n17442), .B1(n7725), .B2(n16942), .ZN(
        n5201) );
  OAI22_X1 U15531 ( .A1(n16945), .A2(n17444), .B1(n7723), .B2(n16942), .ZN(
        n5202) );
  OAI22_X1 U15532 ( .A1(n16945), .A2(n17446), .B1(n7721), .B2(n16942), .ZN(
        n5203) );
  OAI22_X1 U15533 ( .A1(n16945), .A2(n17448), .B1(n7719), .B2(n16942), .ZN(
        n5204) );
  OAI22_X1 U15534 ( .A1(n16945), .A2(n17450), .B1(n7717), .B2(n16942), .ZN(
        n5205) );
  OAI22_X1 U15535 ( .A1(n16946), .A2(n17452), .B1(n7715), .B2(n16942), .ZN(
        n5206) );
  OAI22_X1 U15536 ( .A1(n16946), .A2(n17454), .B1(n7713), .B2(n16942), .ZN(
        n5207) );
  OAI22_X1 U15537 ( .A1(n16946), .A2(n17456), .B1(n7711), .B2(n16943), .ZN(
        n5208) );
  OAI22_X1 U15538 ( .A1(n16946), .A2(n17458), .B1(n7709), .B2(n16943), .ZN(
        n5209) );
  OAI22_X1 U15539 ( .A1(n16946), .A2(n17460), .B1(n7707), .B2(n16943), .ZN(
        n5210) );
  OAI22_X1 U15540 ( .A1(n16947), .A2(n17462), .B1(n7705), .B2(n16943), .ZN(
        n5211) );
  OAI22_X1 U15541 ( .A1(n16947), .A2(n17464), .B1(n7703), .B2(n16943), .ZN(
        n5212) );
  OAI22_X1 U15542 ( .A1(n16947), .A2(n17466), .B1(n7701), .B2(n16943), .ZN(
        n5213) );
  OAI22_X1 U15543 ( .A1(n16947), .A2(n17468), .B1(n7699), .B2(n16943), .ZN(
        n5214) );
  OAI22_X1 U15544 ( .A1(n16947), .A2(n17470), .B1(n7697), .B2(n16943), .ZN(
        n5215) );
  OAI22_X1 U15545 ( .A1(n16948), .A2(n17472), .B1(n7695), .B2(n16943), .ZN(
        n5216) );
  OAI22_X1 U15546 ( .A1(n16948), .A2(n17474), .B1(n7693), .B2(n16943), .ZN(
        n5217) );
  OAI22_X1 U15547 ( .A1(n16948), .A2(n17476), .B1(n7691), .B2(n16943), .ZN(
        n5218) );
  OAI22_X1 U15548 ( .A1(n16948), .A2(n17478), .B1(n7689), .B2(n16943), .ZN(
        n5219) );
  OAI22_X1 U15549 ( .A1(n16995), .A2(n17432), .B1(n7307), .B2(n16993), .ZN(
        n5388) );
  OAI22_X1 U15550 ( .A1(n16995), .A2(n17434), .B1(n7306), .B2(n16993), .ZN(
        n5389) );
  OAI22_X1 U15551 ( .A1(n16995), .A2(n17436), .B1(n7305), .B2(n16993), .ZN(
        n5390) );
  OAI22_X1 U15552 ( .A1(n16995), .A2(n17438), .B1(n7304), .B2(n16993), .ZN(
        n5391) );
  OAI22_X1 U15553 ( .A1(n16995), .A2(n17440), .B1(n7303), .B2(n16993), .ZN(
        n5392) );
  OAI22_X1 U15554 ( .A1(n16996), .A2(n17442), .B1(n7302), .B2(n16993), .ZN(
        n5393) );
  OAI22_X1 U15555 ( .A1(n16996), .A2(n17444), .B1(n7301), .B2(n16993), .ZN(
        n5394) );
  OAI22_X1 U15556 ( .A1(n16996), .A2(n17446), .B1(n7300), .B2(n16993), .ZN(
        n5395) );
  OAI22_X1 U15557 ( .A1(n16996), .A2(n17448), .B1(n7299), .B2(n16993), .ZN(
        n5396) );
  OAI22_X1 U15558 ( .A1(n16996), .A2(n17450), .B1(n7298), .B2(n16993), .ZN(
        n5397) );
  OAI22_X1 U15559 ( .A1(n16997), .A2(n17452), .B1(n7297), .B2(n16993), .ZN(
        n5398) );
  OAI22_X1 U15560 ( .A1(n16997), .A2(n17454), .B1(n7296), .B2(n16993), .ZN(
        n5399) );
  OAI22_X1 U15561 ( .A1(n16997), .A2(n17456), .B1(n7295), .B2(n16994), .ZN(
        n5400) );
  OAI22_X1 U15562 ( .A1(n16997), .A2(n17458), .B1(n7294), .B2(n16994), .ZN(
        n5401) );
  OAI22_X1 U15563 ( .A1(n16997), .A2(n17460), .B1(n7293), .B2(n16994), .ZN(
        n5402) );
  OAI22_X1 U15564 ( .A1(n16998), .A2(n17462), .B1(n7292), .B2(n16994), .ZN(
        n5403) );
  OAI22_X1 U15565 ( .A1(n16998), .A2(n17464), .B1(n7291), .B2(n16994), .ZN(
        n5404) );
  OAI22_X1 U15566 ( .A1(n16998), .A2(n17466), .B1(n7290), .B2(n16994), .ZN(
        n5405) );
  OAI22_X1 U15567 ( .A1(n16998), .A2(n17468), .B1(n7289), .B2(n16994), .ZN(
        n5406) );
  OAI22_X1 U15568 ( .A1(n16998), .A2(n17470), .B1(n7288), .B2(n16994), .ZN(
        n5407) );
  OAI22_X1 U15569 ( .A1(n16999), .A2(n17472), .B1(n7287), .B2(n16994), .ZN(
        n5408) );
  OAI22_X1 U15570 ( .A1(n16999), .A2(n17474), .B1(n7286), .B2(n16994), .ZN(
        n5409) );
  OAI22_X1 U15571 ( .A1(n16999), .A2(n17476), .B1(n7285), .B2(n16994), .ZN(
        n5410) );
  OAI22_X1 U15572 ( .A1(n16999), .A2(n17478), .B1(n7284), .B2(n16994), .ZN(
        n5411) );
  OAI22_X1 U15573 ( .A1(n17012), .A2(n17432), .B1(n8056), .B2(n17010), .ZN(
        n5452) );
  OAI22_X1 U15574 ( .A1(n17012), .A2(n17434), .B1(n8053), .B2(n17010), .ZN(
        n5453) );
  OAI22_X1 U15575 ( .A1(n17012), .A2(n17436), .B1(n8050), .B2(n17010), .ZN(
        n5454) );
  OAI22_X1 U15576 ( .A1(n17012), .A2(n17438), .B1(n8047), .B2(n17010), .ZN(
        n5455) );
  OAI22_X1 U15577 ( .A1(n17012), .A2(n17440), .B1(n8044), .B2(n17010), .ZN(
        n5456) );
  OAI22_X1 U15578 ( .A1(n17013), .A2(n17442), .B1(n8041), .B2(n17010), .ZN(
        n5457) );
  OAI22_X1 U15579 ( .A1(n17013), .A2(n17444), .B1(n8038), .B2(n17010), .ZN(
        n5458) );
  OAI22_X1 U15580 ( .A1(n17013), .A2(n17446), .B1(n8035), .B2(n17010), .ZN(
        n5459) );
  OAI22_X1 U15581 ( .A1(n17013), .A2(n17448), .B1(n8032), .B2(n17010), .ZN(
        n5460) );
  OAI22_X1 U15582 ( .A1(n17013), .A2(n17450), .B1(n8029), .B2(n17010), .ZN(
        n5461) );
  OAI22_X1 U15583 ( .A1(n17014), .A2(n17452), .B1(n8026), .B2(n17010), .ZN(
        n5462) );
  OAI22_X1 U15584 ( .A1(n17014), .A2(n17454), .B1(n8023), .B2(n17010), .ZN(
        n5463) );
  OAI22_X1 U15585 ( .A1(n17014), .A2(n17456), .B1(n8020), .B2(n17011), .ZN(
        n5464) );
  OAI22_X1 U15586 ( .A1(n17014), .A2(n17458), .B1(n8017), .B2(n17011), .ZN(
        n5465) );
  OAI22_X1 U15587 ( .A1(n17014), .A2(n17460), .B1(n8014), .B2(n17011), .ZN(
        n5466) );
  OAI22_X1 U15588 ( .A1(n17015), .A2(n17462), .B1(n8011), .B2(n17011), .ZN(
        n5467) );
  OAI22_X1 U15589 ( .A1(n17015), .A2(n17464), .B1(n8008), .B2(n17011), .ZN(
        n5468) );
  OAI22_X1 U15590 ( .A1(n17015), .A2(n17466), .B1(n8005), .B2(n17011), .ZN(
        n5469) );
  OAI22_X1 U15591 ( .A1(n17015), .A2(n17468), .B1(n8002), .B2(n17011), .ZN(
        n5470) );
  OAI22_X1 U15592 ( .A1(n17015), .A2(n17470), .B1(n7999), .B2(n17011), .ZN(
        n5471) );
  OAI22_X1 U15593 ( .A1(n17016), .A2(n17472), .B1(n7996), .B2(n17011), .ZN(
        n5472) );
  OAI22_X1 U15594 ( .A1(n17016), .A2(n17474), .B1(n7993), .B2(n17011), .ZN(
        n5473) );
  OAI22_X1 U15595 ( .A1(n17016), .A2(n17476), .B1(n7990), .B2(n17011), .ZN(
        n5474) );
  OAI22_X1 U15596 ( .A1(n17016), .A2(n17478), .B1(n7987), .B2(n17011), .ZN(
        n5475) );
  OAI22_X1 U15597 ( .A1(n17029), .A2(n17432), .B1(n8055), .B2(n17027), .ZN(
        n5516) );
  OAI22_X1 U15598 ( .A1(n17029), .A2(n17434), .B1(n8052), .B2(n17027), .ZN(
        n5517) );
  OAI22_X1 U15599 ( .A1(n17029), .A2(n17436), .B1(n8049), .B2(n17027), .ZN(
        n5518) );
  OAI22_X1 U15600 ( .A1(n17029), .A2(n17438), .B1(n8046), .B2(n17027), .ZN(
        n5519) );
  OAI22_X1 U15601 ( .A1(n17029), .A2(n17440), .B1(n8043), .B2(n17027), .ZN(
        n5520) );
  OAI22_X1 U15602 ( .A1(n17030), .A2(n17442), .B1(n8040), .B2(n17027), .ZN(
        n5521) );
  OAI22_X1 U15603 ( .A1(n17030), .A2(n17444), .B1(n8037), .B2(n17027), .ZN(
        n5522) );
  OAI22_X1 U15604 ( .A1(n17030), .A2(n17446), .B1(n8034), .B2(n17027), .ZN(
        n5523) );
  OAI22_X1 U15605 ( .A1(n17030), .A2(n17448), .B1(n8031), .B2(n17027), .ZN(
        n5524) );
  OAI22_X1 U15606 ( .A1(n17030), .A2(n17450), .B1(n8028), .B2(n17027), .ZN(
        n5525) );
  OAI22_X1 U15607 ( .A1(n17031), .A2(n17452), .B1(n8025), .B2(n17027), .ZN(
        n5526) );
  OAI22_X1 U15608 ( .A1(n17031), .A2(n17454), .B1(n8022), .B2(n17027), .ZN(
        n5527) );
  OAI22_X1 U15609 ( .A1(n17031), .A2(n17456), .B1(n8019), .B2(n17028), .ZN(
        n5528) );
  OAI22_X1 U15610 ( .A1(n17031), .A2(n17458), .B1(n8016), .B2(n17028), .ZN(
        n5529) );
  OAI22_X1 U15611 ( .A1(n17031), .A2(n17460), .B1(n8013), .B2(n17028), .ZN(
        n5530) );
  OAI22_X1 U15612 ( .A1(n17032), .A2(n17462), .B1(n8010), .B2(n17028), .ZN(
        n5531) );
  OAI22_X1 U15613 ( .A1(n17032), .A2(n17464), .B1(n8007), .B2(n17028), .ZN(
        n5532) );
  OAI22_X1 U15614 ( .A1(n17032), .A2(n17466), .B1(n8004), .B2(n17028), .ZN(
        n5533) );
  OAI22_X1 U15615 ( .A1(n17032), .A2(n17468), .B1(n8001), .B2(n17028), .ZN(
        n5534) );
  OAI22_X1 U15616 ( .A1(n17032), .A2(n17470), .B1(n7998), .B2(n17028), .ZN(
        n5535) );
  OAI22_X1 U15617 ( .A1(n17033), .A2(n17472), .B1(n7995), .B2(n17028), .ZN(
        n5536) );
  OAI22_X1 U15618 ( .A1(n17033), .A2(n17474), .B1(n7992), .B2(n17028), .ZN(
        n5537) );
  OAI22_X1 U15619 ( .A1(n17033), .A2(n17476), .B1(n7989), .B2(n17028), .ZN(
        n5538) );
  OAI22_X1 U15620 ( .A1(n17033), .A2(n17478), .B1(n7986), .B2(n17028), .ZN(
        n5539) );
  OAI22_X1 U15621 ( .A1(n17046), .A2(n17432), .B1(n7435), .B2(n17044), .ZN(
        n5580) );
  OAI22_X1 U15622 ( .A1(n17046), .A2(n17434), .B1(n7433), .B2(n17044), .ZN(
        n5581) );
  OAI22_X1 U15623 ( .A1(n17046), .A2(n17436), .B1(n7431), .B2(n17044), .ZN(
        n5582) );
  OAI22_X1 U15624 ( .A1(n17046), .A2(n17438), .B1(n7429), .B2(n17044), .ZN(
        n5583) );
  OAI22_X1 U15625 ( .A1(n17046), .A2(n17440), .B1(n7427), .B2(n17044), .ZN(
        n5584) );
  OAI22_X1 U15626 ( .A1(n17047), .A2(n17442), .B1(n7425), .B2(n17044), .ZN(
        n5585) );
  OAI22_X1 U15627 ( .A1(n17047), .A2(n17444), .B1(n7423), .B2(n17044), .ZN(
        n5586) );
  OAI22_X1 U15628 ( .A1(n17047), .A2(n17446), .B1(n7421), .B2(n17044), .ZN(
        n5587) );
  OAI22_X1 U15629 ( .A1(n17047), .A2(n17448), .B1(n7419), .B2(n17044), .ZN(
        n5588) );
  OAI22_X1 U15630 ( .A1(n17047), .A2(n17450), .B1(n7417), .B2(n17044), .ZN(
        n5589) );
  OAI22_X1 U15631 ( .A1(n17048), .A2(n17452), .B1(n7415), .B2(n17044), .ZN(
        n5590) );
  OAI22_X1 U15632 ( .A1(n17048), .A2(n17454), .B1(n7413), .B2(n17044), .ZN(
        n5591) );
  OAI22_X1 U15633 ( .A1(n17048), .A2(n17456), .B1(n7411), .B2(n17045), .ZN(
        n5592) );
  OAI22_X1 U15634 ( .A1(n17048), .A2(n17458), .B1(n7409), .B2(n17045), .ZN(
        n5593) );
  OAI22_X1 U15635 ( .A1(n17048), .A2(n17460), .B1(n7407), .B2(n17045), .ZN(
        n5594) );
  OAI22_X1 U15636 ( .A1(n17049), .A2(n17462), .B1(n7405), .B2(n17045), .ZN(
        n5595) );
  OAI22_X1 U15637 ( .A1(n17049), .A2(n17464), .B1(n7403), .B2(n17045), .ZN(
        n5596) );
  OAI22_X1 U15638 ( .A1(n17049), .A2(n17466), .B1(n7401), .B2(n17045), .ZN(
        n5597) );
  OAI22_X1 U15639 ( .A1(n17049), .A2(n17468), .B1(n7399), .B2(n17045), .ZN(
        n5598) );
  OAI22_X1 U15640 ( .A1(n17049), .A2(n17470), .B1(n7397), .B2(n17045), .ZN(
        n5599) );
  OAI22_X1 U15641 ( .A1(n17050), .A2(n17472), .B1(n7395), .B2(n17045), .ZN(
        n5600) );
  OAI22_X1 U15642 ( .A1(n17050), .A2(n17474), .B1(n7393), .B2(n17045), .ZN(
        n5601) );
  OAI22_X1 U15643 ( .A1(n17050), .A2(n17476), .B1(n7391), .B2(n17045), .ZN(
        n5602) );
  OAI22_X1 U15644 ( .A1(n17050), .A2(n17478), .B1(n7389), .B2(n17045), .ZN(
        n5603) );
  OAI22_X1 U15645 ( .A1(n17173), .A2(n17513), .B1(n988), .B2(n13661), .ZN(
        n6068) );
  OAI22_X1 U15646 ( .A1(n17173), .A2(n17515), .B1(n987), .B2(n17162), .ZN(
        n6069) );
  OAI22_X1 U15647 ( .A1(n17173), .A2(n17517), .B1(n986), .B2(n13661), .ZN(
        n6070) );
  OAI22_X1 U15648 ( .A1(n17173), .A2(n17519), .B1(n985), .B2(n17162), .ZN(
        n6071) );
  OAI22_X1 U15649 ( .A1(n17173), .A2(n17521), .B1(n984), .B2(n13661), .ZN(
        n6072) );
  OAI22_X1 U15650 ( .A1(n17174), .A2(n17523), .B1(n983), .B2(n17162), .ZN(
        n6073) );
  OAI22_X1 U15651 ( .A1(n17174), .A2(n17525), .B1(n982), .B2(n13661), .ZN(
        n6074) );
  OAI22_X1 U15652 ( .A1(n17174), .A2(n17527), .B1(n981), .B2(n17162), .ZN(
        n6075) );
  OAI22_X1 U15653 ( .A1(n17174), .A2(n17529), .B1(n980), .B2(n17163), .ZN(
        n6076) );
  OAI22_X1 U15654 ( .A1(n17174), .A2(n17531), .B1(n979), .B2(n17162), .ZN(
        n6077) );
  OAI22_X1 U15655 ( .A1(n17175), .A2(n17533), .B1(n978), .B2(n17163), .ZN(
        n6078) );
  OAI22_X1 U15656 ( .A1(n17175), .A2(n17535), .B1(n977), .B2(n17162), .ZN(
        n6079) );
  OAI22_X1 U15657 ( .A1(n17175), .A2(n17537), .B1(n976), .B2(n17162), .ZN(
        n6080) );
  OAI22_X1 U15658 ( .A1(n17175), .A2(n17539), .B1(n975), .B2(n17162), .ZN(
        n6081) );
  OAI22_X1 U15659 ( .A1(n17175), .A2(n17541), .B1(n974), .B2(n13661), .ZN(
        n6082) );
  OAI22_X1 U15660 ( .A1(n17176), .A2(n17543), .B1(n973), .B2(n17162), .ZN(
        n6083) );
  OAI22_X1 U15661 ( .A1(n17176), .A2(n17545), .B1(n972), .B2(n13661), .ZN(
        n6084) );
  OAI22_X1 U15662 ( .A1(n17176), .A2(n17547), .B1(n971), .B2(n17162), .ZN(
        n6085) );
  OAI22_X1 U15663 ( .A1(n17176), .A2(n17549), .B1(n970), .B2(n13661), .ZN(
        n6086) );
  OAI22_X1 U15664 ( .A1(n17176), .A2(n17551), .B1(n969), .B2(n17162), .ZN(
        n6087) );
  OAI22_X1 U15665 ( .A1(n17177), .A2(n17553), .B1(n968), .B2(n13661), .ZN(
        n6088) );
  OAI22_X1 U15666 ( .A1(n17177), .A2(n17555), .B1(n967), .B2(n17162), .ZN(
        n6089) );
  OAI22_X1 U15667 ( .A1(n17177), .A2(n17557), .B1(n966), .B2(n13661), .ZN(
        n6090) );
  OAI22_X1 U15668 ( .A1(n17177), .A2(n17578), .B1(n965), .B2(n17162), .ZN(
        n6091) );
  OAI22_X1 U15669 ( .A1(n17183), .A2(n17433), .B1(n964), .B2(n17181), .ZN(
        n6092) );
  OAI22_X1 U15670 ( .A1(n17183), .A2(n17435), .B1(n963), .B2(n17181), .ZN(
        n6093) );
  OAI22_X1 U15671 ( .A1(n17183), .A2(n17437), .B1(n962), .B2(n17181), .ZN(
        n6094) );
  OAI22_X1 U15672 ( .A1(n17183), .A2(n17439), .B1(n961), .B2(n17181), .ZN(
        n6095) );
  OAI22_X1 U15673 ( .A1(n17183), .A2(n17441), .B1(n960), .B2(n17181), .ZN(
        n6096) );
  OAI22_X1 U15674 ( .A1(n17184), .A2(n17443), .B1(n959), .B2(n17181), .ZN(
        n6097) );
  OAI22_X1 U15675 ( .A1(n17184), .A2(n17445), .B1(n958), .B2(n17181), .ZN(
        n6098) );
  OAI22_X1 U15676 ( .A1(n17184), .A2(n17447), .B1(n957), .B2(n17181), .ZN(
        n6099) );
  OAI22_X1 U15677 ( .A1(n17184), .A2(n17449), .B1(n956), .B2(n17181), .ZN(
        n6100) );
  OAI22_X1 U15678 ( .A1(n17184), .A2(n17451), .B1(n955), .B2(n17181), .ZN(
        n6101) );
  OAI22_X1 U15679 ( .A1(n17185), .A2(n17453), .B1(n954), .B2(n17181), .ZN(
        n6102) );
  OAI22_X1 U15680 ( .A1(n17185), .A2(n17455), .B1(n953), .B2(n17181), .ZN(
        n6103) );
  OAI22_X1 U15681 ( .A1(n17185), .A2(n17457), .B1(n952), .B2(n17182), .ZN(
        n6104) );
  OAI22_X1 U15682 ( .A1(n17185), .A2(n17459), .B1(n951), .B2(n17182), .ZN(
        n6105) );
  OAI22_X1 U15683 ( .A1(n17185), .A2(n17461), .B1(n950), .B2(n17182), .ZN(
        n6106) );
  OAI22_X1 U15684 ( .A1(n17186), .A2(n17463), .B1(n949), .B2(n17182), .ZN(
        n6107) );
  OAI22_X1 U15685 ( .A1(n17186), .A2(n17465), .B1(n948), .B2(n17182), .ZN(
        n6108) );
  OAI22_X1 U15686 ( .A1(n17186), .A2(n17467), .B1(n947), .B2(n17182), .ZN(
        n6109) );
  OAI22_X1 U15687 ( .A1(n17186), .A2(n17469), .B1(n946), .B2(n17182), .ZN(
        n6110) );
  OAI22_X1 U15688 ( .A1(n17186), .A2(n17471), .B1(n945), .B2(n17182), .ZN(
        n6111) );
  OAI22_X1 U15689 ( .A1(n17187), .A2(n17473), .B1(n944), .B2(n17182), .ZN(
        n6112) );
  OAI22_X1 U15690 ( .A1(n17187), .A2(n17475), .B1(n943), .B2(n17182), .ZN(
        n6113) );
  OAI22_X1 U15691 ( .A1(n17187), .A2(n17477), .B1(n942), .B2(n17182), .ZN(
        n6114) );
  OAI22_X1 U15692 ( .A1(n17187), .A2(n17479), .B1(n941), .B2(n17182), .ZN(
        n6115) );
  OAI22_X1 U15693 ( .A1(n17322), .A2(n17432), .B1(n16414), .B2(n17319), .ZN(
        n6604) );
  OAI22_X1 U15694 ( .A1(n17322), .A2(n17434), .B1(n16409), .B2(n17319), .ZN(
        n6605) );
  OAI22_X1 U15695 ( .A1(n17322), .A2(n17436), .B1(n16404), .B2(n17319), .ZN(
        n6606) );
  OAI22_X1 U15696 ( .A1(n17322), .A2(n17438), .B1(n16399), .B2(n17319), .ZN(
        n6607) );
  OAI22_X1 U15697 ( .A1(n17322), .A2(n17440), .B1(n16394), .B2(n17319), .ZN(
        n6608) );
  OAI22_X1 U15698 ( .A1(n17323), .A2(n17442), .B1(n16389), .B2(n17319), .ZN(
        n6609) );
  OAI22_X1 U15699 ( .A1(n17323), .A2(n17444), .B1(n16384), .B2(n17319), .ZN(
        n6610) );
  OAI22_X1 U15700 ( .A1(n17323), .A2(n17446), .B1(n16379), .B2(n17319), .ZN(
        n6611) );
  OAI22_X1 U15701 ( .A1(n17323), .A2(n17448), .B1(n16374), .B2(n17319), .ZN(
        n6612) );
  OAI22_X1 U15702 ( .A1(n17323), .A2(n17450), .B1(n16369), .B2(n17319), .ZN(
        n6613) );
  OAI22_X1 U15703 ( .A1(n17324), .A2(n17452), .B1(n16364), .B2(n17319), .ZN(
        n6614) );
  OAI22_X1 U15704 ( .A1(n17324), .A2(n17454), .B1(n16359), .B2(n17319), .ZN(
        n6615) );
  OAI22_X1 U15705 ( .A1(n17324), .A2(n17456), .B1(n16354), .B2(n17320), .ZN(
        n6616) );
  OAI22_X1 U15706 ( .A1(n17324), .A2(n17458), .B1(n16349), .B2(n17320), .ZN(
        n6617) );
  OAI22_X1 U15707 ( .A1(n17324), .A2(n17460), .B1(n16344), .B2(n17320), .ZN(
        n6618) );
  OAI22_X1 U15708 ( .A1(n17325), .A2(n17462), .B1(n16339), .B2(n17320), .ZN(
        n6619) );
  OAI22_X1 U15709 ( .A1(n17325), .A2(n17464), .B1(n16334), .B2(n17320), .ZN(
        n6620) );
  OAI22_X1 U15710 ( .A1(n17325), .A2(n17466), .B1(n16329), .B2(n17320), .ZN(
        n6621) );
  OAI22_X1 U15711 ( .A1(n17325), .A2(n17468), .B1(n16324), .B2(n17320), .ZN(
        n6622) );
  OAI22_X1 U15712 ( .A1(n17325), .A2(n17470), .B1(n16319), .B2(n17320), .ZN(
        n6623) );
  OAI22_X1 U15713 ( .A1(n17326), .A2(n17472), .B1(n16314), .B2(n17320), .ZN(
        n6624) );
  OAI22_X1 U15714 ( .A1(n17326), .A2(n17474), .B1(n16309), .B2(n17320), .ZN(
        n6625) );
  OAI22_X1 U15715 ( .A1(n17326), .A2(n17476), .B1(n16304), .B2(n17320), .ZN(
        n6626) );
  OAI22_X1 U15716 ( .A1(n17326), .A2(n17478), .B1(n16299), .B2(n17320), .ZN(
        n6627) );
  OAI22_X1 U15717 ( .A1(n17341), .A2(n17433), .B1(n7115), .B2(n17338), .ZN(
        n6668) );
  OAI22_X1 U15718 ( .A1(n17341), .A2(n17435), .B1(n7114), .B2(n17338), .ZN(
        n6669) );
  OAI22_X1 U15719 ( .A1(n17341), .A2(n17437), .B1(n7113), .B2(n17338), .ZN(
        n6670) );
  OAI22_X1 U15720 ( .A1(n17341), .A2(n17439), .B1(n7112), .B2(n17338), .ZN(
        n6671) );
  OAI22_X1 U15721 ( .A1(n17341), .A2(n17441), .B1(n7111), .B2(n17338), .ZN(
        n6672) );
  OAI22_X1 U15722 ( .A1(n17342), .A2(n17443), .B1(n7110), .B2(n17338), .ZN(
        n6673) );
  OAI22_X1 U15723 ( .A1(n17342), .A2(n17445), .B1(n7109), .B2(n17338), .ZN(
        n6674) );
  OAI22_X1 U15724 ( .A1(n17342), .A2(n17447), .B1(n7108), .B2(n17338), .ZN(
        n6675) );
  OAI22_X1 U15725 ( .A1(n17342), .A2(n17449), .B1(n7107), .B2(n17338), .ZN(
        n6676) );
  OAI22_X1 U15726 ( .A1(n17342), .A2(n17451), .B1(n7106), .B2(n17338), .ZN(
        n6677) );
  OAI22_X1 U15727 ( .A1(n17343), .A2(n17453), .B1(n7105), .B2(n17338), .ZN(
        n6678) );
  OAI22_X1 U15728 ( .A1(n17343), .A2(n17455), .B1(n7104), .B2(n17338), .ZN(
        n6679) );
  OAI22_X1 U15729 ( .A1(n17343), .A2(n17457), .B1(n7103), .B2(n17339), .ZN(
        n6680) );
  OAI22_X1 U15730 ( .A1(n17343), .A2(n17459), .B1(n7102), .B2(n17339), .ZN(
        n6681) );
  OAI22_X1 U15731 ( .A1(n17343), .A2(n17461), .B1(n7101), .B2(n17339), .ZN(
        n6682) );
  OAI22_X1 U15732 ( .A1(n17344), .A2(n17463), .B1(n7100), .B2(n17339), .ZN(
        n6683) );
  OAI22_X1 U15733 ( .A1(n17344), .A2(n17465), .B1(n7099), .B2(n17339), .ZN(
        n6684) );
  OAI22_X1 U15734 ( .A1(n17344), .A2(n17467), .B1(n7098), .B2(n17339), .ZN(
        n6685) );
  OAI22_X1 U15735 ( .A1(n17344), .A2(n17469), .B1(n7097), .B2(n17339), .ZN(
        n6686) );
  OAI22_X1 U15736 ( .A1(n17344), .A2(n17471), .B1(n7096), .B2(n17339), .ZN(
        n6687) );
  OAI22_X1 U15737 ( .A1(n17345), .A2(n17473), .B1(n7095), .B2(n17339), .ZN(
        n6688) );
  OAI22_X1 U15738 ( .A1(n17345), .A2(n17475), .B1(n7094), .B2(n17339), .ZN(
        n6689) );
  OAI22_X1 U15739 ( .A1(n17345), .A2(n17477), .B1(n7093), .B2(n17339), .ZN(
        n6690) );
  OAI22_X1 U15740 ( .A1(n17345), .A2(n17479), .B1(n7092), .B2(n17339), .ZN(
        n6691) );
  OAI22_X1 U15741 ( .A1(n17360), .A2(n17432), .B1(n16415), .B2(n17357), .ZN(
        n6732) );
  OAI22_X1 U15742 ( .A1(n17360), .A2(n17434), .B1(n16410), .B2(n17357), .ZN(
        n6733) );
  OAI22_X1 U15743 ( .A1(n17360), .A2(n17436), .B1(n16405), .B2(n17357), .ZN(
        n6734) );
  OAI22_X1 U15744 ( .A1(n17360), .A2(n17438), .B1(n16400), .B2(n17357), .ZN(
        n6735) );
  OAI22_X1 U15745 ( .A1(n17360), .A2(n17440), .B1(n16395), .B2(n17357), .ZN(
        n6736) );
  OAI22_X1 U15746 ( .A1(n17361), .A2(n17442), .B1(n16390), .B2(n17357), .ZN(
        n6737) );
  OAI22_X1 U15747 ( .A1(n17361), .A2(n17444), .B1(n16385), .B2(n17357), .ZN(
        n6738) );
  OAI22_X1 U15748 ( .A1(n17361), .A2(n17446), .B1(n16380), .B2(n17357), .ZN(
        n6739) );
  OAI22_X1 U15749 ( .A1(n17361), .A2(n17448), .B1(n16375), .B2(n17357), .ZN(
        n6740) );
  OAI22_X1 U15750 ( .A1(n17361), .A2(n17450), .B1(n16370), .B2(n17357), .ZN(
        n6741) );
  OAI22_X1 U15751 ( .A1(n17362), .A2(n17452), .B1(n16365), .B2(n17357), .ZN(
        n6742) );
  OAI22_X1 U15752 ( .A1(n17362), .A2(n17454), .B1(n16360), .B2(n17357), .ZN(
        n6743) );
  OAI22_X1 U15753 ( .A1(n17362), .A2(n17456), .B1(n16355), .B2(n17358), .ZN(
        n6744) );
  OAI22_X1 U15754 ( .A1(n17362), .A2(n17458), .B1(n16350), .B2(n17358), .ZN(
        n6745) );
  OAI22_X1 U15755 ( .A1(n17362), .A2(n17460), .B1(n16345), .B2(n17358), .ZN(
        n6746) );
  OAI22_X1 U15756 ( .A1(n17363), .A2(n17462), .B1(n16340), .B2(n17358), .ZN(
        n6747) );
  OAI22_X1 U15757 ( .A1(n17363), .A2(n17464), .B1(n16335), .B2(n17358), .ZN(
        n6748) );
  OAI22_X1 U15758 ( .A1(n17363), .A2(n17466), .B1(n16330), .B2(n17358), .ZN(
        n6749) );
  OAI22_X1 U15759 ( .A1(n17363), .A2(n17468), .B1(n16325), .B2(n17358), .ZN(
        n6750) );
  OAI22_X1 U15760 ( .A1(n17363), .A2(n17470), .B1(n16320), .B2(n17358), .ZN(
        n6751) );
  OAI22_X1 U15761 ( .A1(n17364), .A2(n17472), .B1(n16315), .B2(n17358), .ZN(
        n6752) );
  OAI22_X1 U15762 ( .A1(n17364), .A2(n17474), .B1(n16310), .B2(n17358), .ZN(
        n6753) );
  OAI22_X1 U15763 ( .A1(n17364), .A2(n17476), .B1(n16305), .B2(n17358), .ZN(
        n6754) );
  OAI22_X1 U15764 ( .A1(n17364), .A2(n17478), .B1(n16300), .B2(n17358), .ZN(
        n6755) );
  OAI22_X1 U15765 ( .A1(n17379), .A2(n17433), .B1(n16412), .B2(n17376), .ZN(
        n6796) );
  OAI22_X1 U15766 ( .A1(n17379), .A2(n17435), .B1(n16407), .B2(n17376), .ZN(
        n6797) );
  OAI22_X1 U15767 ( .A1(n17379), .A2(n17437), .B1(n16402), .B2(n17376), .ZN(
        n6798) );
  OAI22_X1 U15768 ( .A1(n17379), .A2(n17439), .B1(n16397), .B2(n17376), .ZN(
        n6799) );
  OAI22_X1 U15769 ( .A1(n17379), .A2(n17441), .B1(n16392), .B2(n17376), .ZN(
        n6800) );
  OAI22_X1 U15770 ( .A1(n17380), .A2(n17443), .B1(n16387), .B2(n17376), .ZN(
        n6801) );
  OAI22_X1 U15771 ( .A1(n17380), .A2(n17445), .B1(n16382), .B2(n17376), .ZN(
        n6802) );
  OAI22_X1 U15772 ( .A1(n17380), .A2(n17447), .B1(n16377), .B2(n17376), .ZN(
        n6803) );
  OAI22_X1 U15773 ( .A1(n17380), .A2(n17449), .B1(n16372), .B2(n17376), .ZN(
        n6804) );
  OAI22_X1 U15774 ( .A1(n17380), .A2(n17451), .B1(n16367), .B2(n17376), .ZN(
        n6805) );
  OAI22_X1 U15775 ( .A1(n17381), .A2(n17453), .B1(n16362), .B2(n17376), .ZN(
        n6806) );
  OAI22_X1 U15776 ( .A1(n17381), .A2(n17455), .B1(n16357), .B2(n17376), .ZN(
        n6807) );
  OAI22_X1 U15777 ( .A1(n17381), .A2(n17457), .B1(n16352), .B2(n17377), .ZN(
        n6808) );
  OAI22_X1 U15778 ( .A1(n17381), .A2(n17459), .B1(n16347), .B2(n17377), .ZN(
        n6809) );
  OAI22_X1 U15779 ( .A1(n17381), .A2(n17461), .B1(n16342), .B2(n17377), .ZN(
        n6810) );
  OAI22_X1 U15780 ( .A1(n17382), .A2(n17463), .B1(n16337), .B2(n17377), .ZN(
        n6811) );
  OAI22_X1 U15781 ( .A1(n17382), .A2(n17465), .B1(n16332), .B2(n17377), .ZN(
        n6812) );
  OAI22_X1 U15782 ( .A1(n17382), .A2(n17467), .B1(n16327), .B2(n17377), .ZN(
        n6813) );
  OAI22_X1 U15783 ( .A1(n17382), .A2(n17469), .B1(n16322), .B2(n17377), .ZN(
        n6814) );
  OAI22_X1 U15784 ( .A1(n17382), .A2(n17471), .B1(n16317), .B2(n17377), .ZN(
        n6815) );
  OAI22_X1 U15785 ( .A1(n17383), .A2(n17473), .B1(n16312), .B2(n17377), .ZN(
        n6816) );
  OAI22_X1 U15786 ( .A1(n17383), .A2(n17475), .B1(n16307), .B2(n17377), .ZN(
        n6817) );
  OAI22_X1 U15787 ( .A1(n17383), .A2(n17477), .B1(n16302), .B2(n17377), .ZN(
        n6818) );
  OAI22_X1 U15788 ( .A1(n17383), .A2(n17479), .B1(n16297), .B2(n17377), .ZN(
        n6819) );
  OAI22_X1 U15789 ( .A1(n17417), .A2(n17432), .B1(n8054), .B2(n17414), .ZN(
        n6924) );
  OAI22_X1 U15790 ( .A1(n17417), .A2(n17434), .B1(n8051), .B2(n17414), .ZN(
        n6925) );
  OAI22_X1 U15791 ( .A1(n17417), .A2(n17436), .B1(n8048), .B2(n17414), .ZN(
        n6926) );
  OAI22_X1 U15792 ( .A1(n17417), .A2(n17438), .B1(n8045), .B2(n17414), .ZN(
        n6927) );
  OAI22_X1 U15793 ( .A1(n17417), .A2(n17440), .B1(n8042), .B2(n17414), .ZN(
        n6928) );
  OAI22_X1 U15794 ( .A1(n17418), .A2(n17442), .B1(n8039), .B2(n17414), .ZN(
        n6929) );
  OAI22_X1 U15795 ( .A1(n17418), .A2(n17444), .B1(n8036), .B2(n17414), .ZN(
        n6930) );
  OAI22_X1 U15796 ( .A1(n17418), .A2(n17446), .B1(n8033), .B2(n17414), .ZN(
        n6931) );
  OAI22_X1 U15797 ( .A1(n17418), .A2(n17448), .B1(n8030), .B2(n17414), .ZN(
        n6932) );
  OAI22_X1 U15798 ( .A1(n17418), .A2(n17450), .B1(n8027), .B2(n17414), .ZN(
        n6933) );
  OAI22_X1 U15799 ( .A1(n17419), .A2(n17452), .B1(n8024), .B2(n17414), .ZN(
        n6934) );
  OAI22_X1 U15800 ( .A1(n17419), .A2(n17454), .B1(n8021), .B2(n17414), .ZN(
        n6935) );
  OAI22_X1 U15801 ( .A1(n17419), .A2(n17456), .B1(n8018), .B2(n17415), .ZN(
        n6936) );
  OAI22_X1 U15802 ( .A1(n17419), .A2(n17458), .B1(n8015), .B2(n17415), .ZN(
        n6937) );
  OAI22_X1 U15803 ( .A1(n17419), .A2(n17460), .B1(n8012), .B2(n17415), .ZN(
        n6938) );
  OAI22_X1 U15804 ( .A1(n17420), .A2(n17462), .B1(n8009), .B2(n17415), .ZN(
        n6939) );
  OAI22_X1 U15805 ( .A1(n17420), .A2(n17464), .B1(n8006), .B2(n17415), .ZN(
        n6940) );
  OAI22_X1 U15806 ( .A1(n17420), .A2(n17466), .B1(n8003), .B2(n17415), .ZN(
        n6941) );
  OAI22_X1 U15807 ( .A1(n17420), .A2(n17468), .B1(n8000), .B2(n17415), .ZN(
        n6942) );
  OAI22_X1 U15808 ( .A1(n17420), .A2(n17470), .B1(n7997), .B2(n17415), .ZN(
        n6943) );
  OAI22_X1 U15809 ( .A1(n17421), .A2(n17472), .B1(n7994), .B2(n17415), .ZN(
        n6944) );
  OAI22_X1 U15810 ( .A1(n17421), .A2(n17474), .B1(n7991), .B2(n17415), .ZN(
        n6945) );
  OAI22_X1 U15811 ( .A1(n17421), .A2(n17476), .B1(n7988), .B2(n17415), .ZN(
        n6946) );
  OAI22_X1 U15812 ( .A1(n17421), .A2(n17478), .B1(n7985), .B2(n17415), .ZN(
        n6947) );
  OAI22_X1 U15813 ( .A1(n17562), .A2(n17433), .B1(n7434), .B2(n17559), .ZN(
        n6988) );
  OAI22_X1 U15814 ( .A1(n17562), .A2(n17435), .B1(n7432), .B2(n17559), .ZN(
        n6989) );
  OAI22_X1 U15815 ( .A1(n17562), .A2(n17437), .B1(n7430), .B2(n17559), .ZN(
        n6990) );
  OAI22_X1 U15816 ( .A1(n17562), .A2(n17439), .B1(n7428), .B2(n17559), .ZN(
        n6991) );
  OAI22_X1 U15817 ( .A1(n17562), .A2(n17441), .B1(n7426), .B2(n17559), .ZN(
        n6992) );
  OAI22_X1 U15818 ( .A1(n17563), .A2(n17443), .B1(n7424), .B2(n17559), .ZN(
        n6993) );
  OAI22_X1 U15819 ( .A1(n17563), .A2(n17445), .B1(n7422), .B2(n17559), .ZN(
        n6994) );
  OAI22_X1 U15820 ( .A1(n17563), .A2(n17447), .B1(n7420), .B2(n17559), .ZN(
        n6995) );
  OAI22_X1 U15821 ( .A1(n17563), .A2(n17449), .B1(n7418), .B2(n17559), .ZN(
        n6996) );
  OAI22_X1 U15822 ( .A1(n17563), .A2(n17451), .B1(n7416), .B2(n17559), .ZN(
        n6997) );
  OAI22_X1 U15823 ( .A1(n17564), .A2(n17453), .B1(n7414), .B2(n17559), .ZN(
        n6998) );
  OAI22_X1 U15824 ( .A1(n17564), .A2(n17455), .B1(n7412), .B2(n17559), .ZN(
        n6999) );
  OAI22_X1 U15825 ( .A1(n17564), .A2(n17457), .B1(n7410), .B2(n17560), .ZN(
        n7000) );
  OAI22_X1 U15826 ( .A1(n17564), .A2(n17459), .B1(n7408), .B2(n17560), .ZN(
        n7001) );
  OAI22_X1 U15827 ( .A1(n17564), .A2(n17461), .B1(n7406), .B2(n17560), .ZN(
        n7002) );
  OAI22_X1 U15828 ( .A1(n17565), .A2(n17463), .B1(n7404), .B2(n17560), .ZN(
        n7003) );
  OAI22_X1 U15829 ( .A1(n17565), .A2(n17465), .B1(n7402), .B2(n17560), .ZN(
        n7004) );
  OAI22_X1 U15830 ( .A1(n17565), .A2(n17467), .B1(n7400), .B2(n17560), .ZN(
        n7005) );
  OAI22_X1 U15831 ( .A1(n17565), .A2(n17469), .B1(n7398), .B2(n17560), .ZN(
        n7006) );
  OAI22_X1 U15832 ( .A1(n17565), .A2(n17471), .B1(n7396), .B2(n17560), .ZN(
        n7007) );
  OAI22_X1 U15833 ( .A1(n17566), .A2(n17473), .B1(n7394), .B2(n17560), .ZN(
        n7008) );
  OAI22_X1 U15834 ( .A1(n17566), .A2(n17475), .B1(n7392), .B2(n17560), .ZN(
        n7009) );
  OAI22_X1 U15835 ( .A1(n17566), .A2(n17477), .B1(n7390), .B2(n17560), .ZN(
        n7010) );
  OAI22_X1 U15836 ( .A1(n17566), .A2(n17479), .B1(n7388), .B2(n17560), .ZN(
        n7011) );
  OAI22_X1 U15837 ( .A1(n16931), .A2(n17480), .B1(n7815), .B2(n16925), .ZN(
        n5156) );
  OAI22_X1 U15838 ( .A1(n16932), .A2(n17482), .B1(n7813), .B2(n16926), .ZN(
        n5157) );
  OAI22_X1 U15839 ( .A1(n16932), .A2(n17484), .B1(n7811), .B2(n16924), .ZN(
        n5158) );
  OAI22_X1 U15840 ( .A1(n16932), .A2(n17486), .B1(n7809), .B2(n16925), .ZN(
        n5159) );
  OAI22_X1 U15841 ( .A1(n16932), .A2(n17488), .B1(n7807), .B2(n16926), .ZN(
        n5160) );
  OAI22_X1 U15842 ( .A1(n16932), .A2(n17490), .B1(n7805), .B2(n16924), .ZN(
        n5161) );
  OAI22_X1 U15843 ( .A1(n16933), .A2(n17492), .B1(n7803), .B2(n16925), .ZN(
        n5162) );
  OAI22_X1 U15844 ( .A1(n16933), .A2(n17494), .B1(n7801), .B2(n16926), .ZN(
        n5163) );
  OAI22_X1 U15845 ( .A1(n16933), .A2(n17496), .B1(n7799), .B2(n16924), .ZN(
        n5164) );
  OAI22_X1 U15846 ( .A1(n16933), .A2(n17498), .B1(n7797), .B2(n16925), .ZN(
        n5165) );
  OAI22_X1 U15847 ( .A1(n16933), .A2(n17500), .B1(n7795), .B2(n16926), .ZN(
        n5166) );
  OAI22_X1 U15848 ( .A1(n16934), .A2(n17502), .B1(n7793), .B2(n16924), .ZN(
        n5167) );
  OAI22_X1 U15849 ( .A1(n16934), .A2(n17504), .B1(n7791), .B2(n13677), .ZN(
        n5168) );
  OAI22_X1 U15850 ( .A1(n16934), .A2(n17506), .B1(n7789), .B2(n16924), .ZN(
        n5169) );
  OAI22_X1 U15851 ( .A1(n16934), .A2(n17508), .B1(n7787), .B2(n13677), .ZN(
        n5170) );
  OAI22_X1 U15852 ( .A1(n16934), .A2(n17510), .B1(n7785), .B2(n16924), .ZN(
        n5171) );
  OAI22_X1 U15853 ( .A1(n16935), .A2(n17512), .B1(n7783), .B2(n13677), .ZN(
        n5172) );
  OAI22_X1 U15854 ( .A1(n16935), .A2(n17514), .B1(n7781), .B2(n16924), .ZN(
        n5173) );
  OAI22_X1 U15855 ( .A1(n16935), .A2(n17516), .B1(n7779), .B2(n16925), .ZN(
        n5174) );
  OAI22_X1 U15856 ( .A1(n16935), .A2(n17518), .B1(n7777), .B2(n16926), .ZN(
        n5175) );
  OAI22_X1 U15857 ( .A1(n16935), .A2(n17520), .B1(n7775), .B2(n16924), .ZN(
        n5176) );
  OAI22_X1 U15858 ( .A1(n16936), .A2(n17522), .B1(n7773), .B2(n16924), .ZN(
        n5177) );
  OAI22_X1 U15859 ( .A1(n16936), .A2(n17524), .B1(n7771), .B2(n16925), .ZN(
        n5178) );
  OAI22_X1 U15860 ( .A1(n16936), .A2(n17526), .B1(n7769), .B2(n16926), .ZN(
        n5179) );
  OAI22_X1 U15861 ( .A1(n16936), .A2(n17528), .B1(n7767), .B2(n16924), .ZN(
        n5180) );
  OAI22_X1 U15862 ( .A1(n16936), .A2(n17530), .B1(n7765), .B2(n16924), .ZN(
        n5181) );
  OAI22_X1 U15863 ( .A1(n16937), .A2(n17532), .B1(n7763), .B2(n13677), .ZN(
        n5182) );
  OAI22_X1 U15864 ( .A1(n16937), .A2(n17534), .B1(n7761), .B2(n16924), .ZN(
        n5183) );
  OAI22_X1 U15865 ( .A1(n16937), .A2(n17536), .B1(n7759), .B2(n13677), .ZN(
        n5184) );
  OAI22_X1 U15866 ( .A1(n16937), .A2(n17538), .B1(n7757), .B2(n16924), .ZN(
        n5185) );
  OAI22_X1 U15867 ( .A1(n16937), .A2(n17540), .B1(n7755), .B2(n13677), .ZN(
        n5186) );
  OAI22_X1 U15868 ( .A1(n16938), .A2(n17542), .B1(n7753), .B2(n16924), .ZN(
        n5187) );
  OAI22_X1 U15869 ( .A1(n16938), .A2(n17544), .B1(n7751), .B2(n13677), .ZN(
        n5188) );
  OAI22_X1 U15870 ( .A1(n16938), .A2(n17546), .B1(n7749), .B2(n16924), .ZN(
        n5189) );
  OAI22_X1 U15871 ( .A1(n16938), .A2(n17548), .B1(n7747), .B2(n13677), .ZN(
        n5190) );
  OAI22_X1 U15872 ( .A1(n16938), .A2(n17550), .B1(n7745), .B2(n16924), .ZN(
        n5191) );
  OAI22_X1 U15873 ( .A1(n16948), .A2(n17480), .B1(n7687), .B2(n16942), .ZN(
        n5220) );
  OAI22_X1 U15874 ( .A1(n16949), .A2(n17482), .B1(n7685), .B2(n16943), .ZN(
        n5221) );
  OAI22_X1 U15875 ( .A1(n16949), .A2(n17484), .B1(n7683), .B2(n16941), .ZN(
        n5222) );
  OAI22_X1 U15876 ( .A1(n16949), .A2(n17486), .B1(n7681), .B2(n16942), .ZN(
        n5223) );
  OAI22_X1 U15877 ( .A1(n16949), .A2(n17488), .B1(n7679), .B2(n16943), .ZN(
        n5224) );
  OAI22_X1 U15878 ( .A1(n16949), .A2(n17490), .B1(n7677), .B2(n16941), .ZN(
        n5225) );
  OAI22_X1 U15879 ( .A1(n16950), .A2(n17492), .B1(n7675), .B2(n16942), .ZN(
        n5226) );
  OAI22_X1 U15880 ( .A1(n16950), .A2(n17494), .B1(n7673), .B2(n16943), .ZN(
        n5227) );
  OAI22_X1 U15881 ( .A1(n16950), .A2(n17496), .B1(n7671), .B2(n16941), .ZN(
        n5228) );
  OAI22_X1 U15882 ( .A1(n16950), .A2(n17498), .B1(n7669), .B2(n16942), .ZN(
        n5229) );
  OAI22_X1 U15883 ( .A1(n16950), .A2(n17500), .B1(n7667), .B2(n16943), .ZN(
        n5230) );
  OAI22_X1 U15884 ( .A1(n16951), .A2(n17502), .B1(n7665), .B2(n16941), .ZN(
        n5231) );
  OAI22_X1 U15885 ( .A1(n16951), .A2(n17504), .B1(n7663), .B2(n13676), .ZN(
        n5232) );
  OAI22_X1 U15886 ( .A1(n16951), .A2(n17506), .B1(n7661), .B2(n16941), .ZN(
        n5233) );
  OAI22_X1 U15887 ( .A1(n16951), .A2(n17508), .B1(n7659), .B2(n13676), .ZN(
        n5234) );
  OAI22_X1 U15888 ( .A1(n16951), .A2(n17510), .B1(n7657), .B2(n16941), .ZN(
        n5235) );
  OAI22_X1 U15889 ( .A1(n16952), .A2(n17512), .B1(n7655), .B2(n13676), .ZN(
        n5236) );
  OAI22_X1 U15890 ( .A1(n16952), .A2(n17514), .B1(n7653), .B2(n16941), .ZN(
        n5237) );
  OAI22_X1 U15891 ( .A1(n16952), .A2(n17516), .B1(n7651), .B2(n16942), .ZN(
        n5238) );
  OAI22_X1 U15892 ( .A1(n16952), .A2(n17518), .B1(n7649), .B2(n16943), .ZN(
        n5239) );
  OAI22_X1 U15893 ( .A1(n16952), .A2(n17520), .B1(n7647), .B2(n16941), .ZN(
        n5240) );
  OAI22_X1 U15894 ( .A1(n16953), .A2(n17522), .B1(n7645), .B2(n16941), .ZN(
        n5241) );
  OAI22_X1 U15895 ( .A1(n16953), .A2(n17524), .B1(n7643), .B2(n16942), .ZN(
        n5242) );
  OAI22_X1 U15896 ( .A1(n16953), .A2(n17526), .B1(n7641), .B2(n16943), .ZN(
        n5243) );
  OAI22_X1 U15897 ( .A1(n16953), .A2(n17528), .B1(n7639), .B2(n16941), .ZN(
        n5244) );
  OAI22_X1 U15898 ( .A1(n16953), .A2(n17530), .B1(n7637), .B2(n16941), .ZN(
        n5245) );
  OAI22_X1 U15899 ( .A1(n16954), .A2(n17532), .B1(n7635), .B2(n13676), .ZN(
        n5246) );
  OAI22_X1 U15900 ( .A1(n16954), .A2(n17534), .B1(n7633), .B2(n16941), .ZN(
        n5247) );
  OAI22_X1 U15901 ( .A1(n16954), .A2(n17536), .B1(n7631), .B2(n13676), .ZN(
        n5248) );
  OAI22_X1 U15902 ( .A1(n16954), .A2(n17538), .B1(n7629), .B2(n16941), .ZN(
        n5249) );
  OAI22_X1 U15903 ( .A1(n16954), .A2(n17540), .B1(n7627), .B2(n13676), .ZN(
        n5250) );
  OAI22_X1 U15904 ( .A1(n16955), .A2(n17542), .B1(n7625), .B2(n16941), .ZN(
        n5251) );
  OAI22_X1 U15905 ( .A1(n16955), .A2(n17544), .B1(n7623), .B2(n13676), .ZN(
        n5252) );
  OAI22_X1 U15906 ( .A1(n16955), .A2(n17546), .B1(n7621), .B2(n16941), .ZN(
        n5253) );
  OAI22_X1 U15907 ( .A1(n16955), .A2(n17548), .B1(n7619), .B2(n13676), .ZN(
        n5254) );
  OAI22_X1 U15908 ( .A1(n16955), .A2(n17550), .B1(n7617), .B2(n16941), .ZN(
        n5255) );
  OAI22_X1 U15909 ( .A1(n16999), .A2(n17480), .B1(n7283), .B2(n16993), .ZN(
        n5412) );
  OAI22_X1 U15910 ( .A1(n17000), .A2(n17482), .B1(n7282), .B2(n16994), .ZN(
        n5413) );
  OAI22_X1 U15911 ( .A1(n17000), .A2(n17484), .B1(n7281), .B2(n16992), .ZN(
        n5414) );
  OAI22_X1 U15912 ( .A1(n17000), .A2(n17486), .B1(n7280), .B2(n16993), .ZN(
        n5415) );
  OAI22_X1 U15913 ( .A1(n17000), .A2(n17488), .B1(n7279), .B2(n16994), .ZN(
        n5416) );
  OAI22_X1 U15914 ( .A1(n17000), .A2(n17490), .B1(n7278), .B2(n16992), .ZN(
        n5417) );
  OAI22_X1 U15915 ( .A1(n17001), .A2(n17492), .B1(n7277), .B2(n16993), .ZN(
        n5418) );
  OAI22_X1 U15916 ( .A1(n17001), .A2(n17494), .B1(n7276), .B2(n16994), .ZN(
        n5419) );
  OAI22_X1 U15917 ( .A1(n17001), .A2(n17496), .B1(n7275), .B2(n16992), .ZN(
        n5420) );
  OAI22_X1 U15918 ( .A1(n17001), .A2(n17498), .B1(n7274), .B2(n16993), .ZN(
        n5421) );
  OAI22_X1 U15919 ( .A1(n17001), .A2(n17500), .B1(n7273), .B2(n16994), .ZN(
        n5422) );
  OAI22_X1 U15920 ( .A1(n17002), .A2(n17502), .B1(n7272), .B2(n16992), .ZN(
        n5423) );
  OAI22_X1 U15921 ( .A1(n17002), .A2(n17504), .B1(n7271), .B2(n13673), .ZN(
        n5424) );
  OAI22_X1 U15922 ( .A1(n17002), .A2(n17506), .B1(n7270), .B2(n16992), .ZN(
        n5425) );
  OAI22_X1 U15923 ( .A1(n17002), .A2(n17508), .B1(n7269), .B2(n13673), .ZN(
        n5426) );
  OAI22_X1 U15924 ( .A1(n17002), .A2(n17510), .B1(n7268), .B2(n16992), .ZN(
        n5427) );
  OAI22_X1 U15925 ( .A1(n17003), .A2(n17512), .B1(n7267), .B2(n13673), .ZN(
        n5428) );
  OAI22_X1 U15926 ( .A1(n17003), .A2(n17514), .B1(n7266), .B2(n16992), .ZN(
        n5429) );
  OAI22_X1 U15927 ( .A1(n17003), .A2(n17516), .B1(n7265), .B2(n16993), .ZN(
        n5430) );
  OAI22_X1 U15928 ( .A1(n17003), .A2(n17518), .B1(n7264), .B2(n16994), .ZN(
        n5431) );
  OAI22_X1 U15929 ( .A1(n17003), .A2(n17520), .B1(n7263), .B2(n16992), .ZN(
        n5432) );
  OAI22_X1 U15930 ( .A1(n17004), .A2(n17522), .B1(n7262), .B2(n16992), .ZN(
        n5433) );
  OAI22_X1 U15931 ( .A1(n17004), .A2(n17524), .B1(n7261), .B2(n16993), .ZN(
        n5434) );
  OAI22_X1 U15932 ( .A1(n17004), .A2(n17526), .B1(n7260), .B2(n16994), .ZN(
        n5435) );
  OAI22_X1 U15933 ( .A1(n17004), .A2(n17528), .B1(n7259), .B2(n16992), .ZN(
        n5436) );
  OAI22_X1 U15934 ( .A1(n17004), .A2(n17530), .B1(n7258), .B2(n16992), .ZN(
        n5437) );
  OAI22_X1 U15935 ( .A1(n17005), .A2(n17532), .B1(n7257), .B2(n13673), .ZN(
        n5438) );
  OAI22_X1 U15936 ( .A1(n17005), .A2(n17534), .B1(n7256), .B2(n16992), .ZN(
        n5439) );
  OAI22_X1 U15937 ( .A1(n17005), .A2(n17536), .B1(n7255), .B2(n13673), .ZN(
        n5440) );
  OAI22_X1 U15938 ( .A1(n17005), .A2(n17538), .B1(n7254), .B2(n16992), .ZN(
        n5441) );
  OAI22_X1 U15939 ( .A1(n17005), .A2(n17540), .B1(n7253), .B2(n13673), .ZN(
        n5442) );
  OAI22_X1 U15940 ( .A1(n17006), .A2(n17542), .B1(n7252), .B2(n16992), .ZN(
        n5443) );
  OAI22_X1 U15941 ( .A1(n17006), .A2(n17544), .B1(n7251), .B2(n13673), .ZN(
        n5444) );
  OAI22_X1 U15942 ( .A1(n17006), .A2(n17546), .B1(n7250), .B2(n16992), .ZN(
        n5445) );
  OAI22_X1 U15943 ( .A1(n17006), .A2(n17548), .B1(n7249), .B2(n13673), .ZN(
        n5446) );
  OAI22_X1 U15944 ( .A1(n17006), .A2(n17550), .B1(n7248), .B2(n16992), .ZN(
        n5447) );
  OAI22_X1 U15945 ( .A1(n17016), .A2(n17480), .B1(n7984), .B2(n17010), .ZN(
        n5476) );
  OAI22_X1 U15946 ( .A1(n17017), .A2(n17482), .B1(n7981), .B2(n17011), .ZN(
        n5477) );
  OAI22_X1 U15947 ( .A1(n17017), .A2(n17484), .B1(n7978), .B2(n17009), .ZN(
        n5478) );
  OAI22_X1 U15948 ( .A1(n17017), .A2(n17486), .B1(n7975), .B2(n17010), .ZN(
        n5479) );
  OAI22_X1 U15949 ( .A1(n17017), .A2(n17488), .B1(n7972), .B2(n17011), .ZN(
        n5480) );
  OAI22_X1 U15950 ( .A1(n17017), .A2(n17490), .B1(n7969), .B2(n17009), .ZN(
        n5481) );
  OAI22_X1 U15951 ( .A1(n17018), .A2(n17492), .B1(n7966), .B2(n17010), .ZN(
        n5482) );
  OAI22_X1 U15952 ( .A1(n17018), .A2(n17494), .B1(n7963), .B2(n17011), .ZN(
        n5483) );
  OAI22_X1 U15953 ( .A1(n17018), .A2(n17496), .B1(n7960), .B2(n17009), .ZN(
        n5484) );
  OAI22_X1 U15954 ( .A1(n17018), .A2(n17498), .B1(n7957), .B2(n17010), .ZN(
        n5485) );
  OAI22_X1 U15955 ( .A1(n17018), .A2(n17500), .B1(n7954), .B2(n17011), .ZN(
        n5486) );
  OAI22_X1 U15956 ( .A1(n17019), .A2(n17502), .B1(n7951), .B2(n17009), .ZN(
        n5487) );
  OAI22_X1 U15957 ( .A1(n17019), .A2(n17504), .B1(n7948), .B2(n13671), .ZN(
        n5488) );
  OAI22_X1 U15958 ( .A1(n17019), .A2(n17506), .B1(n7945), .B2(n17009), .ZN(
        n5489) );
  OAI22_X1 U15959 ( .A1(n17019), .A2(n17508), .B1(n7942), .B2(n13671), .ZN(
        n5490) );
  OAI22_X1 U15960 ( .A1(n17019), .A2(n17510), .B1(n7939), .B2(n17009), .ZN(
        n5491) );
  OAI22_X1 U15961 ( .A1(n17020), .A2(n17512), .B1(n7936), .B2(n13671), .ZN(
        n5492) );
  OAI22_X1 U15962 ( .A1(n17020), .A2(n17514), .B1(n7933), .B2(n17009), .ZN(
        n5493) );
  OAI22_X1 U15963 ( .A1(n17020), .A2(n17516), .B1(n7930), .B2(n17010), .ZN(
        n5494) );
  OAI22_X1 U15964 ( .A1(n17020), .A2(n17518), .B1(n7927), .B2(n17011), .ZN(
        n5495) );
  OAI22_X1 U15965 ( .A1(n17020), .A2(n17520), .B1(n7924), .B2(n17009), .ZN(
        n5496) );
  OAI22_X1 U15966 ( .A1(n17021), .A2(n17522), .B1(n7921), .B2(n17009), .ZN(
        n5497) );
  OAI22_X1 U15967 ( .A1(n17021), .A2(n17524), .B1(n7918), .B2(n17010), .ZN(
        n5498) );
  OAI22_X1 U15968 ( .A1(n17021), .A2(n17526), .B1(n7915), .B2(n17011), .ZN(
        n5499) );
  OAI22_X1 U15969 ( .A1(n17021), .A2(n17528), .B1(n7912), .B2(n17009), .ZN(
        n5500) );
  OAI22_X1 U15970 ( .A1(n17021), .A2(n17530), .B1(n7909), .B2(n17009), .ZN(
        n5501) );
  OAI22_X1 U15971 ( .A1(n17022), .A2(n17532), .B1(n7906), .B2(n13671), .ZN(
        n5502) );
  OAI22_X1 U15972 ( .A1(n17022), .A2(n17534), .B1(n7903), .B2(n17009), .ZN(
        n5503) );
  OAI22_X1 U15973 ( .A1(n17022), .A2(n17536), .B1(n7900), .B2(n13671), .ZN(
        n5504) );
  OAI22_X1 U15974 ( .A1(n17022), .A2(n17538), .B1(n7897), .B2(n17009), .ZN(
        n5505) );
  OAI22_X1 U15975 ( .A1(n17022), .A2(n17540), .B1(n7894), .B2(n13671), .ZN(
        n5506) );
  OAI22_X1 U15976 ( .A1(n17023), .A2(n17542), .B1(n7891), .B2(n17009), .ZN(
        n5507) );
  OAI22_X1 U15977 ( .A1(n17023), .A2(n17544), .B1(n7888), .B2(n13671), .ZN(
        n5508) );
  OAI22_X1 U15978 ( .A1(n17023), .A2(n17546), .B1(n7885), .B2(n17009), .ZN(
        n5509) );
  OAI22_X1 U15979 ( .A1(n17023), .A2(n17548), .B1(n7882), .B2(n13671), .ZN(
        n5510) );
  OAI22_X1 U15980 ( .A1(n17023), .A2(n17550), .B1(n7879), .B2(n17009), .ZN(
        n5511) );
  OAI22_X1 U15981 ( .A1(n17033), .A2(n17480), .B1(n7983), .B2(n17027), .ZN(
        n5540) );
  OAI22_X1 U15982 ( .A1(n17034), .A2(n17482), .B1(n7980), .B2(n17028), .ZN(
        n5541) );
  OAI22_X1 U15983 ( .A1(n17034), .A2(n17484), .B1(n7977), .B2(n17026), .ZN(
        n5542) );
  OAI22_X1 U15984 ( .A1(n17034), .A2(n17486), .B1(n7974), .B2(n17027), .ZN(
        n5543) );
  OAI22_X1 U15985 ( .A1(n17034), .A2(n17488), .B1(n7971), .B2(n17028), .ZN(
        n5544) );
  OAI22_X1 U15986 ( .A1(n17034), .A2(n17490), .B1(n7968), .B2(n17026), .ZN(
        n5545) );
  OAI22_X1 U15987 ( .A1(n17035), .A2(n17492), .B1(n7965), .B2(n17027), .ZN(
        n5546) );
  OAI22_X1 U15988 ( .A1(n17035), .A2(n17494), .B1(n7962), .B2(n17028), .ZN(
        n5547) );
  OAI22_X1 U15989 ( .A1(n17035), .A2(n17496), .B1(n7959), .B2(n17026), .ZN(
        n5548) );
  OAI22_X1 U15990 ( .A1(n17035), .A2(n17498), .B1(n7956), .B2(n17027), .ZN(
        n5549) );
  OAI22_X1 U15991 ( .A1(n17035), .A2(n17500), .B1(n7953), .B2(n17028), .ZN(
        n5550) );
  OAI22_X1 U15992 ( .A1(n17036), .A2(n17502), .B1(n7950), .B2(n17026), .ZN(
        n5551) );
  OAI22_X1 U15993 ( .A1(n17036), .A2(n17504), .B1(n7947), .B2(n13670), .ZN(
        n5552) );
  OAI22_X1 U15994 ( .A1(n17036), .A2(n17506), .B1(n7944), .B2(n17026), .ZN(
        n5553) );
  OAI22_X1 U15995 ( .A1(n17036), .A2(n17508), .B1(n7941), .B2(n13670), .ZN(
        n5554) );
  OAI22_X1 U15996 ( .A1(n17036), .A2(n17510), .B1(n7938), .B2(n17026), .ZN(
        n5555) );
  OAI22_X1 U15997 ( .A1(n17037), .A2(n17512), .B1(n7935), .B2(n13670), .ZN(
        n5556) );
  OAI22_X1 U15998 ( .A1(n17037), .A2(n17514), .B1(n7932), .B2(n17026), .ZN(
        n5557) );
  OAI22_X1 U15999 ( .A1(n17037), .A2(n17516), .B1(n7929), .B2(n17027), .ZN(
        n5558) );
  OAI22_X1 U16000 ( .A1(n17037), .A2(n17518), .B1(n7926), .B2(n17028), .ZN(
        n5559) );
  OAI22_X1 U16001 ( .A1(n17037), .A2(n17520), .B1(n7923), .B2(n17026), .ZN(
        n5560) );
  OAI22_X1 U16002 ( .A1(n17038), .A2(n17522), .B1(n7920), .B2(n17026), .ZN(
        n5561) );
  OAI22_X1 U16003 ( .A1(n17038), .A2(n17524), .B1(n7917), .B2(n17027), .ZN(
        n5562) );
  OAI22_X1 U16004 ( .A1(n17038), .A2(n17526), .B1(n7914), .B2(n17028), .ZN(
        n5563) );
  OAI22_X1 U16005 ( .A1(n17038), .A2(n17528), .B1(n7911), .B2(n17026), .ZN(
        n5564) );
  OAI22_X1 U16006 ( .A1(n17038), .A2(n17530), .B1(n7908), .B2(n17026), .ZN(
        n5565) );
  OAI22_X1 U16007 ( .A1(n17039), .A2(n17532), .B1(n7905), .B2(n13670), .ZN(
        n5566) );
  OAI22_X1 U16008 ( .A1(n17039), .A2(n17534), .B1(n7902), .B2(n17026), .ZN(
        n5567) );
  OAI22_X1 U16009 ( .A1(n17039), .A2(n17536), .B1(n7899), .B2(n13670), .ZN(
        n5568) );
  OAI22_X1 U16010 ( .A1(n17039), .A2(n17538), .B1(n7896), .B2(n17026), .ZN(
        n5569) );
  OAI22_X1 U16011 ( .A1(n17039), .A2(n17540), .B1(n7893), .B2(n13670), .ZN(
        n5570) );
  OAI22_X1 U16012 ( .A1(n17040), .A2(n17542), .B1(n7890), .B2(n17026), .ZN(
        n5571) );
  OAI22_X1 U16013 ( .A1(n17040), .A2(n17544), .B1(n7887), .B2(n13670), .ZN(
        n5572) );
  OAI22_X1 U16014 ( .A1(n17040), .A2(n17546), .B1(n7884), .B2(n17026), .ZN(
        n5573) );
  OAI22_X1 U16015 ( .A1(n17040), .A2(n17548), .B1(n7881), .B2(n13670), .ZN(
        n5574) );
  OAI22_X1 U16016 ( .A1(n17040), .A2(n17550), .B1(n7878), .B2(n17026), .ZN(
        n5575) );
  OAI22_X1 U16017 ( .A1(n17050), .A2(n17480), .B1(n7387), .B2(n17044), .ZN(
        n5604) );
  OAI22_X1 U16018 ( .A1(n17051), .A2(n17482), .B1(n7385), .B2(n17045), .ZN(
        n5605) );
  OAI22_X1 U16019 ( .A1(n17051), .A2(n17484), .B1(n7383), .B2(n17043), .ZN(
        n5606) );
  OAI22_X1 U16020 ( .A1(n17051), .A2(n17486), .B1(n7381), .B2(n17044), .ZN(
        n5607) );
  OAI22_X1 U16021 ( .A1(n17051), .A2(n17488), .B1(n7379), .B2(n17045), .ZN(
        n5608) );
  OAI22_X1 U16022 ( .A1(n17051), .A2(n17490), .B1(n7377), .B2(n17043), .ZN(
        n5609) );
  OAI22_X1 U16023 ( .A1(n17052), .A2(n17492), .B1(n7375), .B2(n17044), .ZN(
        n5610) );
  OAI22_X1 U16024 ( .A1(n17052), .A2(n17494), .B1(n7373), .B2(n17045), .ZN(
        n5611) );
  OAI22_X1 U16025 ( .A1(n17052), .A2(n17496), .B1(n7371), .B2(n17043), .ZN(
        n5612) );
  OAI22_X1 U16026 ( .A1(n17052), .A2(n17498), .B1(n7369), .B2(n17044), .ZN(
        n5613) );
  OAI22_X1 U16027 ( .A1(n17052), .A2(n17500), .B1(n7367), .B2(n17045), .ZN(
        n5614) );
  OAI22_X1 U16028 ( .A1(n17053), .A2(n17502), .B1(n7365), .B2(n17043), .ZN(
        n5615) );
  OAI22_X1 U16029 ( .A1(n17053), .A2(n17504), .B1(n7363), .B2(n13669), .ZN(
        n5616) );
  OAI22_X1 U16030 ( .A1(n17053), .A2(n17506), .B1(n7361), .B2(n17043), .ZN(
        n5617) );
  OAI22_X1 U16031 ( .A1(n17053), .A2(n17508), .B1(n7359), .B2(n13669), .ZN(
        n5618) );
  OAI22_X1 U16032 ( .A1(n17053), .A2(n17510), .B1(n7357), .B2(n17043), .ZN(
        n5619) );
  OAI22_X1 U16033 ( .A1(n17054), .A2(n17512), .B1(n7355), .B2(n13669), .ZN(
        n5620) );
  OAI22_X1 U16034 ( .A1(n17054), .A2(n17514), .B1(n7353), .B2(n17043), .ZN(
        n5621) );
  OAI22_X1 U16035 ( .A1(n17054), .A2(n17516), .B1(n7351), .B2(n17044), .ZN(
        n5622) );
  OAI22_X1 U16036 ( .A1(n17054), .A2(n17518), .B1(n7349), .B2(n17045), .ZN(
        n5623) );
  OAI22_X1 U16037 ( .A1(n17054), .A2(n17520), .B1(n7347), .B2(n17043), .ZN(
        n5624) );
  OAI22_X1 U16038 ( .A1(n17055), .A2(n17522), .B1(n7345), .B2(n17043), .ZN(
        n5625) );
  OAI22_X1 U16039 ( .A1(n17055), .A2(n17524), .B1(n7343), .B2(n17044), .ZN(
        n5626) );
  OAI22_X1 U16040 ( .A1(n17055), .A2(n17526), .B1(n7341), .B2(n17045), .ZN(
        n5627) );
  OAI22_X1 U16041 ( .A1(n17055), .A2(n17528), .B1(n7339), .B2(n17043), .ZN(
        n5628) );
  OAI22_X1 U16042 ( .A1(n17055), .A2(n17530), .B1(n7337), .B2(n17043), .ZN(
        n5629) );
  OAI22_X1 U16043 ( .A1(n17056), .A2(n17532), .B1(n7335), .B2(n13669), .ZN(
        n5630) );
  OAI22_X1 U16044 ( .A1(n17056), .A2(n17534), .B1(n7333), .B2(n17043), .ZN(
        n5631) );
  OAI22_X1 U16045 ( .A1(n17056), .A2(n17536), .B1(n7331), .B2(n13669), .ZN(
        n5632) );
  OAI22_X1 U16046 ( .A1(n17056), .A2(n17538), .B1(n7329), .B2(n17043), .ZN(
        n5633) );
  OAI22_X1 U16047 ( .A1(n17056), .A2(n17540), .B1(n7327), .B2(n13669), .ZN(
        n5634) );
  OAI22_X1 U16048 ( .A1(n17057), .A2(n17542), .B1(n7325), .B2(n17043), .ZN(
        n5635) );
  OAI22_X1 U16049 ( .A1(n17057), .A2(n17544), .B1(n7323), .B2(n13669), .ZN(
        n5636) );
  OAI22_X1 U16050 ( .A1(n17057), .A2(n17546), .B1(n7321), .B2(n17043), .ZN(
        n5637) );
  OAI22_X1 U16051 ( .A1(n17057), .A2(n17548), .B1(n7319), .B2(n13669), .ZN(
        n5638) );
  OAI22_X1 U16052 ( .A1(n17057), .A2(n17550), .B1(n7317), .B2(n17043), .ZN(
        n5639) );
  OAI22_X1 U16053 ( .A1(n17187), .A2(n17481), .B1(n940), .B2(n17181), .ZN(
        n6116) );
  OAI22_X1 U16054 ( .A1(n17188), .A2(n17483), .B1(n939), .B2(n17182), .ZN(
        n6117) );
  OAI22_X1 U16055 ( .A1(n17188), .A2(n17485), .B1(n938), .B2(n17180), .ZN(
        n6118) );
  OAI22_X1 U16056 ( .A1(n17188), .A2(n17487), .B1(n937), .B2(n17181), .ZN(
        n6119) );
  OAI22_X1 U16057 ( .A1(n17188), .A2(n17489), .B1(n936), .B2(n17182), .ZN(
        n6120) );
  OAI22_X1 U16058 ( .A1(n17188), .A2(n17491), .B1(n935), .B2(n17180), .ZN(
        n6121) );
  OAI22_X1 U16059 ( .A1(n17189), .A2(n17493), .B1(n934), .B2(n17181), .ZN(
        n6122) );
  OAI22_X1 U16060 ( .A1(n17189), .A2(n17495), .B1(n933), .B2(n17182), .ZN(
        n6123) );
  OAI22_X1 U16061 ( .A1(n17189), .A2(n17497), .B1(n932), .B2(n17180), .ZN(
        n6124) );
  OAI22_X1 U16062 ( .A1(n17189), .A2(n17499), .B1(n931), .B2(n17181), .ZN(
        n6125) );
  OAI22_X1 U16063 ( .A1(n17189), .A2(n17501), .B1(n930), .B2(n17182), .ZN(
        n6126) );
  OAI22_X1 U16064 ( .A1(n17190), .A2(n17503), .B1(n929), .B2(n17180), .ZN(
        n6127) );
  OAI22_X1 U16065 ( .A1(n17190), .A2(n17505), .B1(n928), .B2(n13660), .ZN(
        n6128) );
  OAI22_X1 U16066 ( .A1(n17190), .A2(n17507), .B1(n927), .B2(n17180), .ZN(
        n6129) );
  OAI22_X1 U16067 ( .A1(n17190), .A2(n17509), .B1(n926), .B2(n13660), .ZN(
        n6130) );
  OAI22_X1 U16068 ( .A1(n17190), .A2(n17511), .B1(n925), .B2(n17180), .ZN(
        n6131) );
  OAI22_X1 U16069 ( .A1(n17191), .A2(n17513), .B1(n924), .B2(n13660), .ZN(
        n6132) );
  OAI22_X1 U16070 ( .A1(n17191), .A2(n17515), .B1(n923), .B2(n17180), .ZN(
        n6133) );
  OAI22_X1 U16071 ( .A1(n17191), .A2(n17517), .B1(n922), .B2(n17181), .ZN(
        n6134) );
  OAI22_X1 U16072 ( .A1(n17191), .A2(n17519), .B1(n921), .B2(n17182), .ZN(
        n6135) );
  OAI22_X1 U16073 ( .A1(n17191), .A2(n17521), .B1(n920), .B2(n17180), .ZN(
        n6136) );
  OAI22_X1 U16074 ( .A1(n17192), .A2(n17523), .B1(n919), .B2(n17180), .ZN(
        n6137) );
  OAI22_X1 U16075 ( .A1(n17192), .A2(n17525), .B1(n918), .B2(n17181), .ZN(
        n6138) );
  OAI22_X1 U16076 ( .A1(n17192), .A2(n17527), .B1(n917), .B2(n17182), .ZN(
        n6139) );
  OAI22_X1 U16077 ( .A1(n17192), .A2(n17529), .B1(n916), .B2(n17180), .ZN(
        n6140) );
  OAI22_X1 U16078 ( .A1(n17192), .A2(n17531), .B1(n915), .B2(n17180), .ZN(
        n6141) );
  OAI22_X1 U16079 ( .A1(n17193), .A2(n17533), .B1(n914), .B2(n13660), .ZN(
        n6142) );
  OAI22_X1 U16080 ( .A1(n17193), .A2(n17535), .B1(n913), .B2(n17180), .ZN(
        n6143) );
  OAI22_X1 U16081 ( .A1(n17193), .A2(n17537), .B1(n912), .B2(n13660), .ZN(
        n6144) );
  OAI22_X1 U16082 ( .A1(n17193), .A2(n17539), .B1(n911), .B2(n17180), .ZN(
        n6145) );
  OAI22_X1 U16083 ( .A1(n17193), .A2(n17541), .B1(n910), .B2(n13660), .ZN(
        n6146) );
  OAI22_X1 U16084 ( .A1(n17194), .A2(n17543), .B1(n909), .B2(n17180), .ZN(
        n6147) );
  OAI22_X1 U16085 ( .A1(n17194), .A2(n17545), .B1(n908), .B2(n13660), .ZN(
        n6148) );
  OAI22_X1 U16086 ( .A1(n17194), .A2(n17547), .B1(n907), .B2(n17180), .ZN(
        n6149) );
  OAI22_X1 U16087 ( .A1(n17194), .A2(n17549), .B1(n906), .B2(n13660), .ZN(
        n6150) );
  OAI22_X1 U16088 ( .A1(n17194), .A2(n17551), .B1(n905), .B2(n17180), .ZN(
        n6151) );
  OAI22_X1 U16089 ( .A1(n17326), .A2(n17480), .B1(n16294), .B2(n17321), .ZN(
        n6628) );
  OAI22_X1 U16090 ( .A1(n17327), .A2(n17482), .B1(n16289), .B2(n17321), .ZN(
        n6629) );
  OAI22_X1 U16091 ( .A1(n17327), .A2(n17484), .B1(n16284), .B2(n17321), .ZN(
        n6630) );
  OAI22_X1 U16092 ( .A1(n17327), .A2(n17486), .B1(n16279), .B2(n17321), .ZN(
        n6631) );
  OAI22_X1 U16093 ( .A1(n17327), .A2(n17488), .B1(n16274), .B2(n17321), .ZN(
        n6632) );
  OAI22_X1 U16094 ( .A1(n17327), .A2(n17490), .B1(n16269), .B2(n17321), .ZN(
        n6633) );
  OAI22_X1 U16095 ( .A1(n17328), .A2(n17492), .B1(n16264), .B2(n17321), .ZN(
        n6634) );
  OAI22_X1 U16096 ( .A1(n17328), .A2(n17494), .B1(n16259), .B2(n17321), .ZN(
        n6635) );
  OAI22_X1 U16097 ( .A1(n17328), .A2(n17496), .B1(n16254), .B2(n17321), .ZN(
        n6636) );
  OAI22_X1 U16098 ( .A1(n17328), .A2(n17498), .B1(n16249), .B2(n17321), .ZN(
        n6637) );
  OAI22_X1 U16099 ( .A1(n17328), .A2(n17500), .B1(n16244), .B2(n17321), .ZN(
        n6638) );
  OAI22_X1 U16100 ( .A1(n17329), .A2(n17502), .B1(n16239), .B2(n17321), .ZN(
        n6639) );
  OAI22_X1 U16101 ( .A1(n17329), .A2(n17504), .B1(n16234), .B2(n13648), .ZN(
        n6640) );
  OAI22_X1 U16102 ( .A1(n17329), .A2(n17506), .B1(n16229), .B2(n17318), .ZN(
        n6641) );
  OAI22_X1 U16103 ( .A1(n17329), .A2(n17508), .B1(n16224), .B2(n13648), .ZN(
        n6642) );
  OAI22_X1 U16104 ( .A1(n17329), .A2(n17510), .B1(n16219), .B2(n17318), .ZN(
        n6643) );
  OAI22_X1 U16105 ( .A1(n17330), .A2(n17512), .B1(n16214), .B2(n13648), .ZN(
        n6644) );
  OAI22_X1 U16106 ( .A1(n17330), .A2(n17514), .B1(n16209), .B2(n17318), .ZN(
        n6645) );
  OAI22_X1 U16107 ( .A1(n17330), .A2(n17516), .B1(n16204), .B2(n17319), .ZN(
        n6646) );
  OAI22_X1 U16108 ( .A1(n17330), .A2(n17518), .B1(n16199), .B2(n17320), .ZN(
        n6647) );
  OAI22_X1 U16109 ( .A1(n17330), .A2(n17520), .B1(n16194), .B2(n17321), .ZN(
        n6648) );
  OAI22_X1 U16110 ( .A1(n17331), .A2(n17522), .B1(n16189), .B2(n17318), .ZN(
        n6649) );
  OAI22_X1 U16111 ( .A1(n17331), .A2(n17524), .B1(n16184), .B2(n17319), .ZN(
        n6650) );
  OAI22_X1 U16112 ( .A1(n17331), .A2(n17526), .B1(n16179), .B2(n17320), .ZN(
        n6651) );
  OAI22_X1 U16113 ( .A1(n17331), .A2(n17528), .B1(n16174), .B2(n17318), .ZN(
        n6652) );
  OAI22_X1 U16114 ( .A1(n17331), .A2(n17530), .B1(n16169), .B2(n17318), .ZN(
        n6653) );
  OAI22_X1 U16115 ( .A1(n17332), .A2(n17532), .B1(n16164), .B2(n13648), .ZN(
        n6654) );
  OAI22_X1 U16116 ( .A1(n17332), .A2(n17534), .B1(n16159), .B2(n17318), .ZN(
        n6655) );
  OAI22_X1 U16117 ( .A1(n17332), .A2(n17536), .B1(n16154), .B2(n13648), .ZN(
        n6656) );
  OAI22_X1 U16118 ( .A1(n17332), .A2(n17538), .B1(n16149), .B2(n17318), .ZN(
        n6657) );
  OAI22_X1 U16119 ( .A1(n17332), .A2(n17540), .B1(n16144), .B2(n13648), .ZN(
        n6658) );
  OAI22_X1 U16120 ( .A1(n17333), .A2(n17542), .B1(n16139), .B2(n17318), .ZN(
        n6659) );
  OAI22_X1 U16121 ( .A1(n17333), .A2(n17544), .B1(n16134), .B2(n13648), .ZN(
        n6660) );
  OAI22_X1 U16122 ( .A1(n17333), .A2(n17546), .B1(n16129), .B2(n17318), .ZN(
        n6661) );
  OAI22_X1 U16123 ( .A1(n17333), .A2(n17548), .B1(n16124), .B2(n13648), .ZN(
        n6662) );
  OAI22_X1 U16124 ( .A1(n17333), .A2(n17550), .B1(n16119), .B2(n17318), .ZN(
        n6663) );
  OAI22_X1 U16125 ( .A1(n17345), .A2(n17481), .B1(n7091), .B2(n17340), .ZN(
        n6692) );
  OAI22_X1 U16126 ( .A1(n17346), .A2(n17483), .B1(n7090), .B2(n17340), .ZN(
        n6693) );
  OAI22_X1 U16127 ( .A1(n17346), .A2(n17485), .B1(n7089), .B2(n17340), .ZN(
        n6694) );
  OAI22_X1 U16128 ( .A1(n17346), .A2(n17487), .B1(n7088), .B2(n17340), .ZN(
        n6695) );
  OAI22_X1 U16129 ( .A1(n17346), .A2(n17489), .B1(n7087), .B2(n17340), .ZN(
        n6696) );
  OAI22_X1 U16130 ( .A1(n17346), .A2(n17491), .B1(n7086), .B2(n17340), .ZN(
        n6697) );
  OAI22_X1 U16131 ( .A1(n17347), .A2(n17493), .B1(n7085), .B2(n17340), .ZN(
        n6698) );
  OAI22_X1 U16132 ( .A1(n17347), .A2(n17495), .B1(n7084), .B2(n17340), .ZN(
        n6699) );
  OAI22_X1 U16133 ( .A1(n17347), .A2(n17497), .B1(n7083), .B2(n17340), .ZN(
        n6700) );
  OAI22_X1 U16134 ( .A1(n17347), .A2(n17499), .B1(n7082), .B2(n17340), .ZN(
        n6701) );
  OAI22_X1 U16135 ( .A1(n17347), .A2(n17501), .B1(n7081), .B2(n17340), .ZN(
        n6702) );
  OAI22_X1 U16136 ( .A1(n17348), .A2(n17503), .B1(n7080), .B2(n17340), .ZN(
        n6703) );
  OAI22_X1 U16137 ( .A1(n17348), .A2(n17505), .B1(n7079), .B2(n13646), .ZN(
        n6704) );
  OAI22_X1 U16138 ( .A1(n17348), .A2(n17507), .B1(n7078), .B2(n17337), .ZN(
        n6705) );
  OAI22_X1 U16139 ( .A1(n17348), .A2(n17509), .B1(n7077), .B2(n13646), .ZN(
        n6706) );
  OAI22_X1 U16140 ( .A1(n17348), .A2(n17511), .B1(n7076), .B2(n17337), .ZN(
        n6707) );
  OAI22_X1 U16141 ( .A1(n17349), .A2(n17513), .B1(n7075), .B2(n13646), .ZN(
        n6708) );
  OAI22_X1 U16142 ( .A1(n17349), .A2(n17515), .B1(n7074), .B2(n17337), .ZN(
        n6709) );
  OAI22_X1 U16143 ( .A1(n17349), .A2(n17517), .B1(n7073), .B2(n17338), .ZN(
        n6710) );
  OAI22_X1 U16144 ( .A1(n17349), .A2(n17519), .B1(n7072), .B2(n17339), .ZN(
        n6711) );
  OAI22_X1 U16145 ( .A1(n17349), .A2(n17521), .B1(n7071), .B2(n17340), .ZN(
        n6712) );
  OAI22_X1 U16146 ( .A1(n17350), .A2(n17523), .B1(n7070), .B2(n17337), .ZN(
        n6713) );
  OAI22_X1 U16147 ( .A1(n17350), .A2(n17525), .B1(n7069), .B2(n17338), .ZN(
        n6714) );
  OAI22_X1 U16148 ( .A1(n17350), .A2(n17527), .B1(n7068), .B2(n17339), .ZN(
        n6715) );
  OAI22_X1 U16149 ( .A1(n17350), .A2(n17529), .B1(n7067), .B2(n17337), .ZN(
        n6716) );
  OAI22_X1 U16150 ( .A1(n17350), .A2(n17531), .B1(n7066), .B2(n17337), .ZN(
        n6717) );
  OAI22_X1 U16151 ( .A1(n17351), .A2(n17533), .B1(n7065), .B2(n13646), .ZN(
        n6718) );
  OAI22_X1 U16152 ( .A1(n17351), .A2(n17535), .B1(n7064), .B2(n17337), .ZN(
        n6719) );
  OAI22_X1 U16153 ( .A1(n17351), .A2(n17537), .B1(n7063), .B2(n13646), .ZN(
        n6720) );
  OAI22_X1 U16154 ( .A1(n17351), .A2(n17539), .B1(n7062), .B2(n17337), .ZN(
        n6721) );
  OAI22_X1 U16155 ( .A1(n17351), .A2(n17541), .B1(n7061), .B2(n13646), .ZN(
        n6722) );
  OAI22_X1 U16156 ( .A1(n17352), .A2(n17543), .B1(n7060), .B2(n17337), .ZN(
        n6723) );
  OAI22_X1 U16157 ( .A1(n17352), .A2(n17545), .B1(n7059), .B2(n13646), .ZN(
        n6724) );
  OAI22_X1 U16158 ( .A1(n17352), .A2(n17547), .B1(n7058), .B2(n17337), .ZN(
        n6725) );
  OAI22_X1 U16159 ( .A1(n17352), .A2(n17549), .B1(n7057), .B2(n13646), .ZN(
        n6726) );
  OAI22_X1 U16160 ( .A1(n17352), .A2(n17551), .B1(n7056), .B2(n17337), .ZN(
        n6727) );
  OAI22_X1 U16161 ( .A1(n17364), .A2(n17480), .B1(n16295), .B2(n17359), .ZN(
        n6756) );
  OAI22_X1 U16162 ( .A1(n17365), .A2(n17482), .B1(n16290), .B2(n17359), .ZN(
        n6757) );
  OAI22_X1 U16163 ( .A1(n17365), .A2(n17484), .B1(n16285), .B2(n17359), .ZN(
        n6758) );
  OAI22_X1 U16164 ( .A1(n17365), .A2(n17486), .B1(n16280), .B2(n17359), .ZN(
        n6759) );
  OAI22_X1 U16165 ( .A1(n17365), .A2(n17488), .B1(n16275), .B2(n17359), .ZN(
        n6760) );
  OAI22_X1 U16166 ( .A1(n17365), .A2(n17490), .B1(n16270), .B2(n17359), .ZN(
        n6761) );
  OAI22_X1 U16167 ( .A1(n17366), .A2(n17492), .B1(n16265), .B2(n17359), .ZN(
        n6762) );
  OAI22_X1 U16168 ( .A1(n17366), .A2(n17494), .B1(n16260), .B2(n17359), .ZN(
        n6763) );
  OAI22_X1 U16169 ( .A1(n17366), .A2(n17496), .B1(n16255), .B2(n17359), .ZN(
        n6764) );
  OAI22_X1 U16170 ( .A1(n17366), .A2(n17498), .B1(n16250), .B2(n17359), .ZN(
        n6765) );
  OAI22_X1 U16171 ( .A1(n17366), .A2(n17500), .B1(n16245), .B2(n17359), .ZN(
        n6766) );
  OAI22_X1 U16172 ( .A1(n17367), .A2(n17502), .B1(n16240), .B2(n17359), .ZN(
        n6767) );
  OAI22_X1 U16173 ( .A1(n17367), .A2(n17504), .B1(n16235), .B2(n13644), .ZN(
        n6768) );
  OAI22_X1 U16174 ( .A1(n17367), .A2(n17506), .B1(n16230), .B2(n17356), .ZN(
        n6769) );
  OAI22_X1 U16175 ( .A1(n17367), .A2(n17508), .B1(n16225), .B2(n13644), .ZN(
        n6770) );
  OAI22_X1 U16176 ( .A1(n17367), .A2(n17510), .B1(n16220), .B2(n17356), .ZN(
        n6771) );
  OAI22_X1 U16177 ( .A1(n17368), .A2(n17512), .B1(n16215), .B2(n13644), .ZN(
        n6772) );
  OAI22_X1 U16178 ( .A1(n17368), .A2(n17514), .B1(n16210), .B2(n17356), .ZN(
        n6773) );
  OAI22_X1 U16179 ( .A1(n17368), .A2(n17516), .B1(n16205), .B2(n17357), .ZN(
        n6774) );
  OAI22_X1 U16180 ( .A1(n17368), .A2(n17518), .B1(n16200), .B2(n17358), .ZN(
        n6775) );
  OAI22_X1 U16181 ( .A1(n17368), .A2(n17520), .B1(n16195), .B2(n17359), .ZN(
        n6776) );
  OAI22_X1 U16182 ( .A1(n17369), .A2(n17522), .B1(n16190), .B2(n17356), .ZN(
        n6777) );
  OAI22_X1 U16183 ( .A1(n17369), .A2(n17524), .B1(n16185), .B2(n17357), .ZN(
        n6778) );
  OAI22_X1 U16184 ( .A1(n17369), .A2(n17526), .B1(n16180), .B2(n17358), .ZN(
        n6779) );
  OAI22_X1 U16185 ( .A1(n17369), .A2(n17528), .B1(n16175), .B2(n17356), .ZN(
        n6780) );
  OAI22_X1 U16186 ( .A1(n17369), .A2(n17530), .B1(n16170), .B2(n17356), .ZN(
        n6781) );
  OAI22_X1 U16187 ( .A1(n17370), .A2(n17532), .B1(n16165), .B2(n13644), .ZN(
        n6782) );
  OAI22_X1 U16188 ( .A1(n17370), .A2(n17534), .B1(n16160), .B2(n17356), .ZN(
        n6783) );
  OAI22_X1 U16189 ( .A1(n17370), .A2(n17536), .B1(n16155), .B2(n13644), .ZN(
        n6784) );
  OAI22_X1 U16190 ( .A1(n17370), .A2(n17538), .B1(n16150), .B2(n17356), .ZN(
        n6785) );
  OAI22_X1 U16191 ( .A1(n17370), .A2(n17540), .B1(n16145), .B2(n13644), .ZN(
        n6786) );
  OAI22_X1 U16192 ( .A1(n17371), .A2(n17542), .B1(n16140), .B2(n17356), .ZN(
        n6787) );
  OAI22_X1 U16193 ( .A1(n17371), .A2(n17544), .B1(n16135), .B2(n13644), .ZN(
        n6788) );
  OAI22_X1 U16194 ( .A1(n17371), .A2(n17546), .B1(n16130), .B2(n17356), .ZN(
        n6789) );
  OAI22_X1 U16195 ( .A1(n17371), .A2(n17548), .B1(n16125), .B2(n13644), .ZN(
        n6790) );
  OAI22_X1 U16196 ( .A1(n17371), .A2(n17550), .B1(n16120), .B2(n17356), .ZN(
        n6791) );
  OAI22_X1 U16197 ( .A1(n17383), .A2(n17481), .B1(n16292), .B2(n17378), .ZN(
        n6820) );
  OAI22_X1 U16198 ( .A1(n17384), .A2(n17483), .B1(n16287), .B2(n17378), .ZN(
        n6821) );
  OAI22_X1 U16199 ( .A1(n17384), .A2(n17485), .B1(n16282), .B2(n17378), .ZN(
        n6822) );
  OAI22_X1 U16200 ( .A1(n17384), .A2(n17487), .B1(n16277), .B2(n17378), .ZN(
        n6823) );
  OAI22_X1 U16201 ( .A1(n17384), .A2(n17489), .B1(n16272), .B2(n17378), .ZN(
        n6824) );
  OAI22_X1 U16202 ( .A1(n17384), .A2(n17491), .B1(n16267), .B2(n17378), .ZN(
        n6825) );
  OAI22_X1 U16203 ( .A1(n17385), .A2(n17493), .B1(n16262), .B2(n17378), .ZN(
        n6826) );
  OAI22_X1 U16204 ( .A1(n17385), .A2(n17495), .B1(n16257), .B2(n17378), .ZN(
        n6827) );
  OAI22_X1 U16205 ( .A1(n17385), .A2(n17497), .B1(n16252), .B2(n17378), .ZN(
        n6828) );
  OAI22_X1 U16206 ( .A1(n17385), .A2(n17499), .B1(n16247), .B2(n17378), .ZN(
        n6829) );
  OAI22_X1 U16207 ( .A1(n17385), .A2(n17501), .B1(n16242), .B2(n17378), .ZN(
        n6830) );
  OAI22_X1 U16208 ( .A1(n17386), .A2(n17503), .B1(n16237), .B2(n17378), .ZN(
        n6831) );
  OAI22_X1 U16209 ( .A1(n17386), .A2(n17505), .B1(n16232), .B2(n13642), .ZN(
        n6832) );
  OAI22_X1 U16210 ( .A1(n17386), .A2(n17507), .B1(n16227), .B2(n17375), .ZN(
        n6833) );
  OAI22_X1 U16211 ( .A1(n17386), .A2(n17509), .B1(n16222), .B2(n13642), .ZN(
        n6834) );
  OAI22_X1 U16212 ( .A1(n17386), .A2(n17511), .B1(n16217), .B2(n17375), .ZN(
        n6835) );
  OAI22_X1 U16213 ( .A1(n17387), .A2(n17513), .B1(n16212), .B2(n13642), .ZN(
        n6836) );
  OAI22_X1 U16214 ( .A1(n17387), .A2(n17515), .B1(n16207), .B2(n17375), .ZN(
        n6837) );
  OAI22_X1 U16215 ( .A1(n17387), .A2(n17517), .B1(n16202), .B2(n17376), .ZN(
        n6838) );
  OAI22_X1 U16216 ( .A1(n17387), .A2(n17519), .B1(n16197), .B2(n17377), .ZN(
        n6839) );
  OAI22_X1 U16217 ( .A1(n17387), .A2(n17521), .B1(n16192), .B2(n17378), .ZN(
        n6840) );
  OAI22_X1 U16218 ( .A1(n17388), .A2(n17523), .B1(n16187), .B2(n17375), .ZN(
        n6841) );
  OAI22_X1 U16219 ( .A1(n17388), .A2(n17525), .B1(n16182), .B2(n17376), .ZN(
        n6842) );
  OAI22_X1 U16220 ( .A1(n17388), .A2(n17527), .B1(n16177), .B2(n17377), .ZN(
        n6843) );
  OAI22_X1 U16221 ( .A1(n17388), .A2(n17529), .B1(n16172), .B2(n17375), .ZN(
        n6844) );
  OAI22_X1 U16222 ( .A1(n17388), .A2(n17531), .B1(n16167), .B2(n17375), .ZN(
        n6845) );
  OAI22_X1 U16223 ( .A1(n17389), .A2(n17533), .B1(n16162), .B2(n13642), .ZN(
        n6846) );
  OAI22_X1 U16224 ( .A1(n17389), .A2(n17535), .B1(n16157), .B2(n17375), .ZN(
        n6847) );
  OAI22_X1 U16225 ( .A1(n17389), .A2(n17537), .B1(n16152), .B2(n13642), .ZN(
        n6848) );
  OAI22_X1 U16226 ( .A1(n17389), .A2(n17539), .B1(n16147), .B2(n17375), .ZN(
        n6849) );
  OAI22_X1 U16227 ( .A1(n17389), .A2(n17541), .B1(n16142), .B2(n13642), .ZN(
        n6850) );
  OAI22_X1 U16228 ( .A1(n17390), .A2(n17543), .B1(n16137), .B2(n17375), .ZN(
        n6851) );
  OAI22_X1 U16229 ( .A1(n17390), .A2(n17545), .B1(n16132), .B2(n13642), .ZN(
        n6852) );
  OAI22_X1 U16230 ( .A1(n17390), .A2(n17547), .B1(n16127), .B2(n17375), .ZN(
        n6853) );
  OAI22_X1 U16231 ( .A1(n17390), .A2(n17549), .B1(n16122), .B2(n13642), .ZN(
        n6854) );
  OAI22_X1 U16232 ( .A1(n17390), .A2(n17551), .B1(n16117), .B2(n17375), .ZN(
        n6855) );
  OAI22_X1 U16233 ( .A1(n17421), .A2(n17480), .B1(n7982), .B2(n17416), .ZN(
        n6948) );
  OAI22_X1 U16234 ( .A1(n17422), .A2(n17482), .B1(n7979), .B2(n17416), .ZN(
        n6949) );
  OAI22_X1 U16235 ( .A1(n17422), .A2(n17484), .B1(n7976), .B2(n17416), .ZN(
        n6950) );
  OAI22_X1 U16236 ( .A1(n17422), .A2(n17486), .B1(n7973), .B2(n17416), .ZN(
        n6951) );
  OAI22_X1 U16237 ( .A1(n17422), .A2(n17488), .B1(n7970), .B2(n17416), .ZN(
        n6952) );
  OAI22_X1 U16238 ( .A1(n17422), .A2(n17490), .B1(n7967), .B2(n17416), .ZN(
        n6953) );
  OAI22_X1 U16239 ( .A1(n17423), .A2(n17492), .B1(n7964), .B2(n17416), .ZN(
        n6954) );
  OAI22_X1 U16240 ( .A1(n17423), .A2(n17494), .B1(n7961), .B2(n17416), .ZN(
        n6955) );
  OAI22_X1 U16241 ( .A1(n17423), .A2(n17496), .B1(n7958), .B2(n17416), .ZN(
        n6956) );
  OAI22_X1 U16242 ( .A1(n17423), .A2(n17498), .B1(n7955), .B2(n17416), .ZN(
        n6957) );
  OAI22_X1 U16243 ( .A1(n17423), .A2(n17500), .B1(n7952), .B2(n17416), .ZN(
        n6958) );
  OAI22_X1 U16244 ( .A1(n17424), .A2(n17502), .B1(n7949), .B2(n17416), .ZN(
        n6959) );
  OAI22_X1 U16245 ( .A1(n17424), .A2(n17504), .B1(n7946), .B2(n13638), .ZN(
        n6960) );
  OAI22_X1 U16246 ( .A1(n17424), .A2(n17506), .B1(n7943), .B2(n17413), .ZN(
        n6961) );
  OAI22_X1 U16247 ( .A1(n17424), .A2(n17508), .B1(n7940), .B2(n13638), .ZN(
        n6962) );
  OAI22_X1 U16248 ( .A1(n17424), .A2(n17510), .B1(n7937), .B2(n17413), .ZN(
        n6963) );
  OAI22_X1 U16249 ( .A1(n17425), .A2(n17512), .B1(n7934), .B2(n13638), .ZN(
        n6964) );
  OAI22_X1 U16250 ( .A1(n17425), .A2(n17514), .B1(n7931), .B2(n17413), .ZN(
        n6965) );
  OAI22_X1 U16251 ( .A1(n17425), .A2(n17516), .B1(n7928), .B2(n17414), .ZN(
        n6966) );
  OAI22_X1 U16252 ( .A1(n17425), .A2(n17518), .B1(n7925), .B2(n17415), .ZN(
        n6967) );
  OAI22_X1 U16253 ( .A1(n17425), .A2(n17520), .B1(n7922), .B2(n17416), .ZN(
        n6968) );
  OAI22_X1 U16254 ( .A1(n17426), .A2(n17522), .B1(n7919), .B2(n17413), .ZN(
        n6969) );
  OAI22_X1 U16255 ( .A1(n17426), .A2(n17524), .B1(n7916), .B2(n17414), .ZN(
        n6970) );
  OAI22_X1 U16256 ( .A1(n17426), .A2(n17526), .B1(n7913), .B2(n17415), .ZN(
        n6971) );
  OAI22_X1 U16257 ( .A1(n17426), .A2(n17528), .B1(n7910), .B2(n17413), .ZN(
        n6972) );
  OAI22_X1 U16258 ( .A1(n17426), .A2(n17530), .B1(n7907), .B2(n17413), .ZN(
        n6973) );
  OAI22_X1 U16259 ( .A1(n17427), .A2(n17532), .B1(n7904), .B2(n13638), .ZN(
        n6974) );
  OAI22_X1 U16260 ( .A1(n17427), .A2(n17534), .B1(n7901), .B2(n17413), .ZN(
        n6975) );
  OAI22_X1 U16261 ( .A1(n17427), .A2(n17536), .B1(n7898), .B2(n13638), .ZN(
        n6976) );
  OAI22_X1 U16262 ( .A1(n17427), .A2(n17538), .B1(n7895), .B2(n17413), .ZN(
        n6977) );
  OAI22_X1 U16263 ( .A1(n17427), .A2(n17540), .B1(n7892), .B2(n13638), .ZN(
        n6978) );
  OAI22_X1 U16264 ( .A1(n17428), .A2(n17542), .B1(n7889), .B2(n17413), .ZN(
        n6979) );
  OAI22_X1 U16265 ( .A1(n17428), .A2(n17544), .B1(n7886), .B2(n13638), .ZN(
        n6980) );
  OAI22_X1 U16266 ( .A1(n17428), .A2(n17546), .B1(n7883), .B2(n17413), .ZN(
        n6981) );
  OAI22_X1 U16267 ( .A1(n17428), .A2(n17548), .B1(n7880), .B2(n13638), .ZN(
        n6982) );
  OAI22_X1 U16268 ( .A1(n17428), .A2(n17550), .B1(n7877), .B2(n17413), .ZN(
        n6983) );
  OAI22_X1 U16269 ( .A1(n17566), .A2(n17481), .B1(n7386), .B2(n17561), .ZN(
        n7012) );
  OAI22_X1 U16270 ( .A1(n17567), .A2(n17483), .B1(n7384), .B2(n17561), .ZN(
        n7013) );
  OAI22_X1 U16271 ( .A1(n17567), .A2(n17485), .B1(n7382), .B2(n17561), .ZN(
        n7014) );
  OAI22_X1 U16272 ( .A1(n17567), .A2(n17487), .B1(n7380), .B2(n17561), .ZN(
        n7015) );
  OAI22_X1 U16273 ( .A1(n17567), .A2(n17489), .B1(n7378), .B2(n17561), .ZN(
        n7016) );
  OAI22_X1 U16274 ( .A1(n17567), .A2(n17491), .B1(n7376), .B2(n17561), .ZN(
        n7017) );
  OAI22_X1 U16275 ( .A1(n17568), .A2(n17493), .B1(n7374), .B2(n17561), .ZN(
        n7018) );
  OAI22_X1 U16276 ( .A1(n17568), .A2(n17495), .B1(n7372), .B2(n17561), .ZN(
        n7019) );
  OAI22_X1 U16277 ( .A1(n17568), .A2(n17497), .B1(n7370), .B2(n17561), .ZN(
        n7020) );
  OAI22_X1 U16278 ( .A1(n17568), .A2(n17499), .B1(n7368), .B2(n17561), .ZN(
        n7021) );
  OAI22_X1 U16279 ( .A1(n17568), .A2(n17501), .B1(n7366), .B2(n17561), .ZN(
        n7022) );
  OAI22_X1 U16280 ( .A1(n17569), .A2(n17503), .B1(n7364), .B2(n17561), .ZN(
        n7023) );
  OAI22_X1 U16281 ( .A1(n17569), .A2(n17505), .B1(n7362), .B2(n13572), .ZN(
        n7024) );
  OAI22_X1 U16282 ( .A1(n17569), .A2(n17507), .B1(n7360), .B2(n17558), .ZN(
        n7025) );
  OAI22_X1 U16283 ( .A1(n17569), .A2(n17509), .B1(n7358), .B2(n13572), .ZN(
        n7026) );
  OAI22_X1 U16284 ( .A1(n17569), .A2(n17511), .B1(n7356), .B2(n17558), .ZN(
        n7027) );
  OAI22_X1 U16285 ( .A1(n17570), .A2(n17513), .B1(n7354), .B2(n13572), .ZN(
        n7028) );
  OAI22_X1 U16286 ( .A1(n17570), .A2(n17515), .B1(n7352), .B2(n17558), .ZN(
        n7029) );
  OAI22_X1 U16287 ( .A1(n17570), .A2(n17517), .B1(n7350), .B2(n17559), .ZN(
        n7030) );
  OAI22_X1 U16288 ( .A1(n17570), .A2(n17519), .B1(n7348), .B2(n17560), .ZN(
        n7031) );
  OAI22_X1 U16289 ( .A1(n17570), .A2(n17521), .B1(n7346), .B2(n17561), .ZN(
        n7032) );
  OAI22_X1 U16290 ( .A1(n17571), .A2(n17523), .B1(n7344), .B2(n17558), .ZN(
        n7033) );
  OAI22_X1 U16291 ( .A1(n17571), .A2(n17525), .B1(n7342), .B2(n17559), .ZN(
        n7034) );
  OAI22_X1 U16292 ( .A1(n17571), .A2(n17527), .B1(n7340), .B2(n17560), .ZN(
        n7035) );
  OAI22_X1 U16293 ( .A1(n17571), .A2(n17529), .B1(n7338), .B2(n17558), .ZN(
        n7036) );
  OAI22_X1 U16294 ( .A1(n17571), .A2(n17531), .B1(n7336), .B2(n17558), .ZN(
        n7037) );
  OAI22_X1 U16295 ( .A1(n17572), .A2(n17533), .B1(n7334), .B2(n13572), .ZN(
        n7038) );
  OAI22_X1 U16296 ( .A1(n17572), .A2(n17535), .B1(n7332), .B2(n17558), .ZN(
        n7039) );
  OAI22_X1 U16297 ( .A1(n17572), .A2(n17537), .B1(n7330), .B2(n13572), .ZN(
        n7040) );
  OAI22_X1 U16298 ( .A1(n17572), .A2(n17539), .B1(n7328), .B2(n17558), .ZN(
        n7041) );
  OAI22_X1 U16299 ( .A1(n17572), .A2(n17541), .B1(n7326), .B2(n13572), .ZN(
        n7042) );
  OAI22_X1 U16300 ( .A1(n17573), .A2(n17543), .B1(n7324), .B2(n17558), .ZN(
        n7043) );
  OAI22_X1 U16301 ( .A1(n17573), .A2(n17545), .B1(n7322), .B2(n13572), .ZN(
        n7044) );
  OAI22_X1 U16302 ( .A1(n17573), .A2(n17547), .B1(n7320), .B2(n17558), .ZN(
        n7045) );
  OAI22_X1 U16303 ( .A1(n17573), .A2(n17549), .B1(n7318), .B2(n13572), .ZN(
        n7046) );
  OAI22_X1 U16304 ( .A1(n17573), .A2(n17551), .B1(n7316), .B2(n17558), .ZN(
        n7047) );
  OAI22_X1 U16305 ( .A1(n17170), .A2(n17491), .B1(n999), .B2(n17163), .ZN(
        n6057) );
  OAI22_X1 U16306 ( .A1(n17171), .A2(n17493), .B1(n998), .B2(n17163), .ZN(
        n6058) );
  OAI22_X1 U16307 ( .A1(n17171), .A2(n17495), .B1(n997), .B2(n17163), .ZN(
        n6059) );
  OAI22_X1 U16308 ( .A1(n17171), .A2(n17497), .B1(n996), .B2(n17163), .ZN(
        n6060) );
  OAI22_X1 U16309 ( .A1(n17171), .A2(n17499), .B1(n995), .B2(n17163), .ZN(
        n6061) );
  OAI22_X1 U16310 ( .A1(n17171), .A2(n17501), .B1(n994), .B2(n17163), .ZN(
        n6062) );
  OAI22_X1 U16311 ( .A1(n17172), .A2(n17503), .B1(n993), .B2(n17163), .ZN(
        n6063) );
  OAI22_X1 U16312 ( .A1(n17172), .A2(n17505), .B1(n992), .B2(n17163), .ZN(
        n6064) );
  OAI22_X1 U16313 ( .A1(n17172), .A2(n17507), .B1(n991), .B2(n17163), .ZN(
        n6065) );
  OAI22_X1 U16314 ( .A1(n17172), .A2(n17509), .B1(n990), .B2(n17163), .ZN(
        n6066) );
  OAI22_X1 U16315 ( .A1(n17172), .A2(n17511), .B1(n989), .B2(n17163), .ZN(
        n6067) );
  OAI22_X1 U16316 ( .A1(n16939), .A2(n17552), .B1(n7743), .B2(n13677), .ZN(
        n5192) );
  OAI22_X1 U16317 ( .A1(n16939), .A2(n17554), .B1(n7741), .B2(n13677), .ZN(
        n5193) );
  OAI22_X1 U16318 ( .A1(n16939), .A2(n17556), .B1(n7739), .B2(n16924), .ZN(
        n5194) );
  OAI22_X1 U16319 ( .A1(n16939), .A2(n17577), .B1(n7737), .B2(n13677), .ZN(
        n5195) );
  OAI22_X1 U16320 ( .A1(n17041), .A2(n17552), .B1(n7875), .B2(n13670), .ZN(
        n5576) );
  OAI22_X1 U16321 ( .A1(n17041), .A2(n17554), .B1(n7872), .B2(n13670), .ZN(
        n5577) );
  OAI22_X1 U16322 ( .A1(n17041), .A2(n17556), .B1(n7869), .B2(n17026), .ZN(
        n5578) );
  OAI22_X1 U16323 ( .A1(n17041), .A2(n17577), .B1(n7866), .B2(n13670), .ZN(
        n5579) );
  OAI22_X1 U16324 ( .A1(n17195), .A2(n17553), .B1(n904), .B2(n13660), .ZN(
        n6152) );
  OAI22_X1 U16325 ( .A1(n17195), .A2(n17555), .B1(n903), .B2(n13660), .ZN(
        n6153) );
  OAI22_X1 U16326 ( .A1(n17195), .A2(n17557), .B1(n902), .B2(n17180), .ZN(
        n6154) );
  OAI22_X1 U16327 ( .A1(n17195), .A2(n17578), .B1(n901), .B2(n13660), .ZN(
        n6155) );
  OAI22_X1 U16328 ( .A1(n17334), .A2(n17552), .B1(n16114), .B2(n13648), .ZN(
        n6664) );
  OAI22_X1 U16329 ( .A1(n17334), .A2(n17554), .B1(n16109), .B2(n13648), .ZN(
        n6665) );
  OAI22_X1 U16330 ( .A1(n17334), .A2(n17556), .B1(n16104), .B2(n17318), .ZN(
        n6666) );
  OAI22_X1 U16331 ( .A1(n17334), .A2(n17577), .B1(n16099), .B2(n13648), .ZN(
        n6667) );
  OAI22_X1 U16332 ( .A1(n17391), .A2(n17553), .B1(n16112), .B2(n13642), .ZN(
        n6856) );
  OAI22_X1 U16333 ( .A1(n17391), .A2(n17555), .B1(n16107), .B2(n13642), .ZN(
        n6857) );
  OAI22_X1 U16334 ( .A1(n17391), .A2(n17557), .B1(n16102), .B2(n17375), .ZN(
        n6858) );
  OAI22_X1 U16335 ( .A1(n17391), .A2(n17578), .B1(n16097), .B2(n13642), .ZN(
        n6859) );
  OAI22_X1 U16336 ( .A1(n16956), .A2(n17552), .B1(n7615), .B2(n13676), .ZN(
        n5256) );
  OAI22_X1 U16337 ( .A1(n16956), .A2(n17554), .B1(n7613), .B2(n13676), .ZN(
        n5257) );
  OAI22_X1 U16338 ( .A1(n16956), .A2(n17556), .B1(n7611), .B2(n16941), .ZN(
        n5258) );
  OAI22_X1 U16339 ( .A1(n16956), .A2(n17577), .B1(n7609), .B2(n13676), .ZN(
        n5259) );
  OAI22_X1 U16340 ( .A1(n17007), .A2(n17552), .B1(n7247), .B2(n13673), .ZN(
        n5448) );
  OAI22_X1 U16341 ( .A1(n17007), .A2(n17554), .B1(n7246), .B2(n13673), .ZN(
        n5449) );
  OAI22_X1 U16342 ( .A1(n17007), .A2(n17556), .B1(n7245), .B2(n16992), .ZN(
        n5450) );
  OAI22_X1 U16343 ( .A1(n17007), .A2(n17577), .B1(n7244), .B2(n13673), .ZN(
        n5451) );
  OAI22_X1 U16344 ( .A1(n17024), .A2(n17552), .B1(n7876), .B2(n13671), .ZN(
        n5512) );
  OAI22_X1 U16345 ( .A1(n17024), .A2(n17554), .B1(n7873), .B2(n13671), .ZN(
        n5513) );
  OAI22_X1 U16346 ( .A1(n17024), .A2(n17556), .B1(n7870), .B2(n17009), .ZN(
        n5514) );
  OAI22_X1 U16347 ( .A1(n17024), .A2(n17577), .B1(n7867), .B2(n13671), .ZN(
        n5515) );
  OAI22_X1 U16348 ( .A1(n17058), .A2(n17552), .B1(n7315), .B2(n13669), .ZN(
        n5640) );
  OAI22_X1 U16349 ( .A1(n17058), .A2(n17554), .B1(n7313), .B2(n13669), .ZN(
        n5641) );
  OAI22_X1 U16350 ( .A1(n17058), .A2(n17556), .B1(n7311), .B2(n17043), .ZN(
        n5642) );
  OAI22_X1 U16351 ( .A1(n17058), .A2(n17577), .B1(n7309), .B2(n13669), .ZN(
        n5643) );
  OAI22_X1 U16352 ( .A1(n17353), .A2(n17552), .B1(n7055), .B2(n13646), .ZN(
        n6728) );
  OAI22_X1 U16353 ( .A1(n17353), .A2(n17554), .B1(n7054), .B2(n13646), .ZN(
        n6729) );
  OAI22_X1 U16354 ( .A1(n17353), .A2(n17556), .B1(n7053), .B2(n17337), .ZN(
        n6730) );
  OAI22_X1 U16355 ( .A1(n17353), .A2(n17577), .B1(n7052), .B2(n13646), .ZN(
        n6731) );
  OAI22_X1 U16356 ( .A1(n17372), .A2(n17553), .B1(n16115), .B2(n13644), .ZN(
        n6792) );
  OAI22_X1 U16357 ( .A1(n17372), .A2(n17555), .B1(n16110), .B2(n13644), .ZN(
        n6793) );
  OAI22_X1 U16358 ( .A1(n17372), .A2(n17557), .B1(n16105), .B2(n17356), .ZN(
        n6794) );
  OAI22_X1 U16359 ( .A1(n17372), .A2(n17578), .B1(n16100), .B2(n13644), .ZN(
        n6795) );
  OAI22_X1 U16360 ( .A1(n17429), .A2(n17552), .B1(n7874), .B2(n13638), .ZN(
        n6984) );
  OAI22_X1 U16361 ( .A1(n17429), .A2(n17554), .B1(n7871), .B2(n13638), .ZN(
        n6985) );
  OAI22_X1 U16362 ( .A1(n17429), .A2(n17556), .B1(n7868), .B2(n17413), .ZN(
        n6986) );
  OAI22_X1 U16363 ( .A1(n17429), .A2(n17577), .B1(n7865), .B2(n13638), .ZN(
        n6987) );
  OAI22_X1 U16364 ( .A1(n17574), .A2(n17553), .B1(n7314), .B2(n13572), .ZN(
        n7048) );
  OAI22_X1 U16365 ( .A1(n17574), .A2(n17555), .B1(n7312), .B2(n13572), .ZN(
        n7049) );
  OAI22_X1 U16366 ( .A1(n17574), .A2(n17557), .B1(n7310), .B2(n17558), .ZN(
        n7050) );
  OAI22_X1 U16367 ( .A1(n17574), .A2(n17578), .B1(n7308), .B2(n13572), .ZN(
        n7051) );
  OAI22_X1 U16368 ( .A1(n16973), .A2(n17552), .B1(n13675), .B2(n13318), .ZN(
        n5320) );
  OAI22_X1 U16369 ( .A1(n16973), .A2(n17554), .B1(n13675), .B2(n13317), .ZN(
        n5321) );
  OAI22_X1 U16370 ( .A1(n16973), .A2(n17556), .B1(n16958), .B2(n13316), .ZN(
        n5322) );
  OAI22_X1 U16371 ( .A1(n16973), .A2(n17577), .B1(n13675), .B2(n13315), .ZN(
        n5323) );
  OAI22_X1 U16372 ( .A1(n16990), .A2(n17552), .B1(n13674), .B2(n13254), .ZN(
        n5384) );
  OAI22_X1 U16373 ( .A1(n16990), .A2(n17554), .B1(n13674), .B2(n13253), .ZN(
        n5385) );
  OAI22_X1 U16374 ( .A1(n16990), .A2(n17556), .B1(n16975), .B2(n13252), .ZN(
        n5386) );
  OAI22_X1 U16375 ( .A1(n16990), .A2(n17577), .B1(n13674), .B2(n13251), .ZN(
        n5387) );
  OAI22_X1 U16376 ( .A1(n17092), .A2(n17552), .B1(n13667), .B2(n12934), .ZN(
        n5768) );
  OAI22_X1 U16377 ( .A1(n17092), .A2(n17554), .B1(n13667), .B2(n12933), .ZN(
        n5769) );
  OAI22_X1 U16378 ( .A1(n17092), .A2(n17556), .B1(n17077), .B2(n12932), .ZN(
        n5770) );
  OAI22_X1 U16379 ( .A1(n17092), .A2(n17577), .B1(n13667), .B2(n12931), .ZN(
        n5771) );
  OAI22_X1 U16380 ( .A1(n17143), .A2(n17553), .B1(n13664), .B2(n12870), .ZN(
        n5960) );
  OAI22_X1 U16381 ( .A1(n17143), .A2(n17555), .B1(n13664), .B2(n12869), .ZN(
        n5961) );
  OAI22_X1 U16382 ( .A1(n17143), .A2(n17557), .B1(n17128), .B2(n12868), .ZN(
        n5962) );
  OAI22_X1 U16383 ( .A1(n17143), .A2(n17578), .B1(n13664), .B2(n12867), .ZN(
        n5963) );
  OAI22_X1 U16384 ( .A1(n17160), .A2(n17553), .B1(n13662), .B2(n12806), .ZN(
        n6024) );
  OAI22_X1 U16385 ( .A1(n17160), .A2(n17555), .B1(n13662), .B2(n12805), .ZN(
        n6025) );
  OAI22_X1 U16386 ( .A1(n17160), .A2(n17557), .B1(n17145), .B2(n12804), .ZN(
        n6026) );
  OAI22_X1 U16387 ( .A1(n17160), .A2(n17578), .B1(n13662), .B2(n12803), .ZN(
        n6027) );
  OAI22_X1 U16388 ( .A1(n17246), .A2(n17553), .B1(n13657), .B2(n12649), .ZN(
        n6344) );
  OAI22_X1 U16389 ( .A1(n17246), .A2(n17555), .B1(n13657), .B2(n12648), .ZN(
        n6345) );
  OAI22_X1 U16390 ( .A1(n17246), .A2(n17557), .B1(n17231), .B2(n12647), .ZN(
        n6346) );
  OAI22_X1 U16391 ( .A1(n17246), .A2(n17578), .B1(n13657), .B2(n12646), .ZN(
        n6347) );
  OAI22_X1 U16392 ( .A1(n17280), .A2(n17553), .B1(n13655), .B2(n12521), .ZN(
        n6472) );
  OAI22_X1 U16393 ( .A1(n17280), .A2(n17555), .B1(n13655), .B2(n12520), .ZN(
        n6473) );
  OAI22_X1 U16394 ( .A1(n17280), .A2(n17557), .B1(n17265), .B2(n12519), .ZN(
        n6474) );
  OAI22_X1 U16395 ( .A1(n17280), .A2(n17578), .B1(n13655), .B2(n12518), .ZN(
        n6475) );
  OAI22_X1 U16396 ( .A1(n17297), .A2(n17553), .B1(n13653), .B2(n12457), .ZN(
        n6536) );
  OAI22_X1 U16397 ( .A1(n17297), .A2(n17555), .B1(n13653), .B2(n12456), .ZN(
        n6537) );
  OAI22_X1 U16398 ( .A1(n17297), .A2(n17557), .B1(n17282), .B2(n12455), .ZN(
        n6538) );
  OAI22_X1 U16399 ( .A1(n17297), .A2(n17578), .B1(n13653), .B2(n12454), .ZN(
        n6539) );
  NAND2_X1 U16400 ( .A1(n16056), .A2(n16057), .ZN(n4876) );
  NOR4_X1 U16401 ( .A1(n16077), .A2(n16078), .A3(n16079), .A4(n16080), .ZN(
        n16056) );
  NOR4_X1 U16402 ( .A1(n16058), .A2(n16059), .A3(n16060), .A4(n16061), .ZN(
        n16057) );
  OAI221_X1 U16403 ( .B1(n16411), .B2(n16554), .C1(n16412), .C2(n16548), .A(
        n16084), .ZN(n16079) );
  NAND2_X1 U16404 ( .A1(n15534), .A2(n15535), .ZN(n4905) );
  NOR4_X1 U16405 ( .A1(n15544), .A2(n15545), .A3(n15546), .A4(n15547), .ZN(
        n15534) );
  NOR4_X1 U16406 ( .A1(n15536), .A2(n15537), .A3(n15538), .A4(n15539), .ZN(
        n15535) );
  OAI221_X1 U16407 ( .B1(n13477), .B2(n16532), .C1(n999), .C2(n16526), .A(
        n15550), .ZN(n15545) );
  NAND2_X1 U16408 ( .A1(n15516), .A2(n15517), .ZN(n4906) );
  NOR4_X1 U16409 ( .A1(n15526), .A2(n15527), .A3(n15528), .A4(n15529), .ZN(
        n15516) );
  NOR4_X1 U16410 ( .A1(n15518), .A2(n15519), .A3(n15520), .A4(n15521), .ZN(
        n15517) );
  OAI221_X1 U16411 ( .B1(n13476), .B2(n16532), .C1(n998), .C2(n16526), .A(
        n15532), .ZN(n15527) );
  NAND2_X1 U16412 ( .A1(n15498), .A2(n15499), .ZN(n4907) );
  NOR4_X1 U16413 ( .A1(n15508), .A2(n15509), .A3(n15510), .A4(n15511), .ZN(
        n15498) );
  NOR4_X1 U16414 ( .A1(n15500), .A2(n15501), .A3(n15502), .A4(n15503), .ZN(
        n15499) );
  OAI221_X1 U16415 ( .B1(n13475), .B2(n16532), .C1(n997), .C2(n16526), .A(
        n15514), .ZN(n15509) );
  NAND2_X1 U16416 ( .A1(n15480), .A2(n15481), .ZN(n4908) );
  NOR4_X1 U16417 ( .A1(n15490), .A2(n15491), .A3(n15492), .A4(n15493), .ZN(
        n15480) );
  NOR4_X1 U16418 ( .A1(n15482), .A2(n15483), .A3(n15484), .A4(n15485), .ZN(
        n15481) );
  OAI221_X1 U16419 ( .B1(n13474), .B2(n16532), .C1(n996), .C2(n16526), .A(
        n15496), .ZN(n15491) );
  NAND2_X1 U16420 ( .A1(n15462), .A2(n15463), .ZN(n4909) );
  NOR4_X1 U16421 ( .A1(n15472), .A2(n15473), .A3(n15474), .A4(n15475), .ZN(
        n15462) );
  NOR4_X1 U16422 ( .A1(n15464), .A2(n15465), .A3(n15466), .A4(n15467), .ZN(
        n15463) );
  OAI221_X1 U16423 ( .B1(n13473), .B2(n16532), .C1(n995), .C2(n16526), .A(
        n15478), .ZN(n15473) );
  NAND2_X1 U16424 ( .A1(n15444), .A2(n15445), .ZN(n4910) );
  NOR4_X1 U16425 ( .A1(n15454), .A2(n15455), .A3(n15456), .A4(n15457), .ZN(
        n15444) );
  NOR4_X1 U16426 ( .A1(n15446), .A2(n15447), .A3(n15448), .A4(n15449), .ZN(
        n15445) );
  OAI221_X1 U16427 ( .B1(n13472), .B2(n16532), .C1(n994), .C2(n16526), .A(
        n15460), .ZN(n15455) );
  NAND2_X1 U16428 ( .A1(n15426), .A2(n15427), .ZN(n4911) );
  NOR4_X1 U16429 ( .A1(n15436), .A2(n15437), .A3(n15438), .A4(n15439), .ZN(
        n15426) );
  NOR4_X1 U16430 ( .A1(n15428), .A2(n15429), .A3(n15430), .A4(n15431), .ZN(
        n15427) );
  OAI221_X1 U16431 ( .B1(n13471), .B2(n16532), .C1(n993), .C2(n16526), .A(
        n15442), .ZN(n15437) );
  NAND2_X1 U16432 ( .A1(n15408), .A2(n15409), .ZN(n4912) );
  NOR4_X1 U16433 ( .A1(n15418), .A2(n15419), .A3(n15420), .A4(n15421), .ZN(
        n15408) );
  NOR4_X1 U16434 ( .A1(n15410), .A2(n15411), .A3(n15412), .A4(n15413), .ZN(
        n15409) );
  OAI221_X1 U16435 ( .B1(n13470), .B2(n16533), .C1(n992), .C2(n16527), .A(
        n15424), .ZN(n15419) );
  NAND2_X1 U16436 ( .A1(n15390), .A2(n15391), .ZN(n4913) );
  NOR4_X1 U16437 ( .A1(n15400), .A2(n15401), .A3(n15402), .A4(n15403), .ZN(
        n15390) );
  NOR4_X1 U16438 ( .A1(n15392), .A2(n15393), .A3(n15394), .A4(n15395), .ZN(
        n15391) );
  OAI221_X1 U16439 ( .B1(n13469), .B2(n16533), .C1(n991), .C2(n16527), .A(
        n15406), .ZN(n15401) );
  NAND2_X1 U16440 ( .A1(n15372), .A2(n15373), .ZN(n4914) );
  NOR4_X1 U16441 ( .A1(n15382), .A2(n15383), .A3(n15384), .A4(n15385), .ZN(
        n15372) );
  NOR4_X1 U16442 ( .A1(n15374), .A2(n15375), .A3(n15376), .A4(n15377), .ZN(
        n15373) );
  OAI221_X1 U16443 ( .B1(n13468), .B2(n16533), .C1(n990), .C2(n16527), .A(
        n15388), .ZN(n15383) );
  NAND2_X1 U16444 ( .A1(n15354), .A2(n15355), .ZN(n4915) );
  NOR4_X1 U16445 ( .A1(n15364), .A2(n15365), .A3(n15366), .A4(n15367), .ZN(
        n15354) );
  NOR4_X1 U16446 ( .A1(n15356), .A2(n15357), .A3(n15358), .A4(n15359), .ZN(
        n15355) );
  OAI221_X1 U16447 ( .B1(n13467), .B2(n16533), .C1(n989), .C2(n16527), .A(
        n15370), .ZN(n15365) );
  NAND2_X1 U16448 ( .A1(n15336), .A2(n15337), .ZN(n4916) );
  NOR4_X1 U16449 ( .A1(n15346), .A2(n15347), .A3(n15348), .A4(n15349), .ZN(
        n15336) );
  NOR4_X1 U16450 ( .A1(n15338), .A2(n15339), .A3(n15340), .A4(n15341), .ZN(
        n15337) );
  OAI221_X1 U16451 ( .B1(n13466), .B2(n16533), .C1(n988), .C2(n16527), .A(
        n15352), .ZN(n15347) );
  NAND2_X1 U16452 ( .A1(n15318), .A2(n15319), .ZN(n4917) );
  NOR4_X1 U16453 ( .A1(n15328), .A2(n15329), .A3(n15330), .A4(n15331), .ZN(
        n15318) );
  NOR4_X1 U16454 ( .A1(n15320), .A2(n15321), .A3(n15322), .A4(n15323), .ZN(
        n15319) );
  OAI221_X1 U16455 ( .B1(n13465), .B2(n16533), .C1(n987), .C2(n16527), .A(
        n15334), .ZN(n15329) );
  NAND2_X1 U16456 ( .A1(n15300), .A2(n15301), .ZN(n4918) );
  NOR4_X1 U16457 ( .A1(n15310), .A2(n15311), .A3(n15312), .A4(n15313), .ZN(
        n15300) );
  NOR4_X1 U16458 ( .A1(n15302), .A2(n15303), .A3(n15304), .A4(n15305), .ZN(
        n15301) );
  OAI221_X1 U16459 ( .B1(n13464), .B2(n16533), .C1(n986), .C2(n16527), .A(
        n15316), .ZN(n15311) );
  NAND2_X1 U16460 ( .A1(n15282), .A2(n15283), .ZN(n4919) );
  NOR4_X1 U16461 ( .A1(n15292), .A2(n15293), .A3(n15294), .A4(n15295), .ZN(
        n15282) );
  NOR4_X1 U16462 ( .A1(n15284), .A2(n15285), .A3(n15286), .A4(n15287), .ZN(
        n15283) );
  OAI221_X1 U16463 ( .B1(n13463), .B2(n16533), .C1(n985), .C2(n16527), .A(
        n15298), .ZN(n15293) );
  NAND2_X1 U16464 ( .A1(n15264), .A2(n15265), .ZN(n4920) );
  NOR4_X1 U16465 ( .A1(n15274), .A2(n15275), .A3(n15276), .A4(n15277), .ZN(
        n15264) );
  NOR4_X1 U16466 ( .A1(n15266), .A2(n15267), .A3(n15268), .A4(n15269), .ZN(
        n15265) );
  OAI221_X1 U16467 ( .B1(n13462), .B2(n16533), .C1(n984), .C2(n16527), .A(
        n15280), .ZN(n15275) );
  NAND2_X1 U16468 ( .A1(n15246), .A2(n15247), .ZN(n4921) );
  NOR4_X1 U16469 ( .A1(n15256), .A2(n15257), .A3(n15258), .A4(n15259), .ZN(
        n15246) );
  NOR4_X1 U16470 ( .A1(n15248), .A2(n15249), .A3(n15250), .A4(n15251), .ZN(
        n15247) );
  OAI221_X1 U16471 ( .B1(n13461), .B2(n16533), .C1(n983), .C2(n16527), .A(
        n15262), .ZN(n15257) );
  NAND2_X1 U16472 ( .A1(n15228), .A2(n15229), .ZN(n4922) );
  NOR4_X1 U16473 ( .A1(n15238), .A2(n15239), .A3(n15240), .A4(n15241), .ZN(
        n15228) );
  NOR4_X1 U16474 ( .A1(n15230), .A2(n15231), .A3(n15232), .A4(n15233), .ZN(
        n15229) );
  OAI221_X1 U16475 ( .B1(n13460), .B2(n16533), .C1(n982), .C2(n16527), .A(
        n15244), .ZN(n15239) );
  NAND2_X1 U16476 ( .A1(n15210), .A2(n15211), .ZN(n4923) );
  NOR4_X1 U16477 ( .A1(n15220), .A2(n15221), .A3(n15222), .A4(n15223), .ZN(
        n15210) );
  NOR4_X1 U16478 ( .A1(n15212), .A2(n15213), .A3(n15214), .A4(n15215), .ZN(
        n15211) );
  OAI221_X1 U16479 ( .B1(n13459), .B2(n16533), .C1(n981), .C2(n16527), .A(
        n15226), .ZN(n15221) );
  NAND2_X1 U16480 ( .A1(n14848), .A2(n14849), .ZN(n4940) );
  NOR4_X1 U16481 ( .A1(n14869), .A2(n14870), .A3(n14871), .A4(n14872), .ZN(
        n14848) );
  NOR4_X1 U16482 ( .A1(n14850), .A2(n14851), .A3(n14852), .A4(n14853), .ZN(
        n14849) );
  OAI221_X1 U16483 ( .B1(n16411), .B2(n16759), .C1(n16412), .C2(n16753), .A(
        n14876), .ZN(n14871) );
  NAND2_X1 U16484 ( .A1(n14830), .A2(n14831), .ZN(n4941) );
  NOR4_X1 U16485 ( .A1(n14840), .A2(n14841), .A3(n14842), .A4(n14843), .ZN(
        n14830) );
  NOR4_X1 U16486 ( .A1(n14832), .A2(n14833), .A3(n14834), .A4(n14835), .ZN(
        n14831) );
  OAI221_X1 U16487 ( .B1(n16406), .B2(n16759), .C1(n16407), .C2(n16753), .A(
        n14845), .ZN(n14842) );
  NAND2_X1 U16488 ( .A1(n14812), .A2(n14813), .ZN(n4942) );
  NOR4_X1 U16489 ( .A1(n14822), .A2(n14823), .A3(n14824), .A4(n14825), .ZN(
        n14812) );
  NOR4_X1 U16490 ( .A1(n14814), .A2(n14815), .A3(n14816), .A4(n14817), .ZN(
        n14813) );
  OAI221_X1 U16491 ( .B1(n16401), .B2(n16759), .C1(n16402), .C2(n16753), .A(
        n14827), .ZN(n14824) );
  NAND2_X1 U16492 ( .A1(n14794), .A2(n14795), .ZN(n4943) );
  NOR4_X1 U16493 ( .A1(n14804), .A2(n14805), .A3(n14806), .A4(n14807), .ZN(
        n14794) );
  NOR4_X1 U16494 ( .A1(n14796), .A2(n14797), .A3(n14798), .A4(n14799), .ZN(
        n14795) );
  OAI221_X1 U16495 ( .B1(n16396), .B2(n16759), .C1(n16397), .C2(n16753), .A(
        n14809), .ZN(n14806) );
  NAND2_X1 U16496 ( .A1(n14776), .A2(n14777), .ZN(n4944) );
  NOR4_X1 U16497 ( .A1(n14786), .A2(n14787), .A3(n14788), .A4(n14789), .ZN(
        n14776) );
  NOR4_X1 U16498 ( .A1(n14778), .A2(n14779), .A3(n14780), .A4(n14781), .ZN(
        n14777) );
  OAI221_X1 U16499 ( .B1(n16391), .B2(n16759), .C1(n16392), .C2(n16753), .A(
        n14791), .ZN(n14788) );
  NAND2_X1 U16500 ( .A1(n14758), .A2(n14759), .ZN(n4945) );
  NOR4_X1 U16501 ( .A1(n14768), .A2(n14769), .A3(n14770), .A4(n14771), .ZN(
        n14758) );
  NOR4_X1 U16502 ( .A1(n14760), .A2(n14761), .A3(n14762), .A4(n14763), .ZN(
        n14759) );
  OAI221_X1 U16503 ( .B1(n16386), .B2(n16759), .C1(n16387), .C2(n16753), .A(
        n14773), .ZN(n14770) );
  NAND2_X1 U16504 ( .A1(n14740), .A2(n14741), .ZN(n4946) );
  NOR4_X1 U16505 ( .A1(n14750), .A2(n14751), .A3(n14752), .A4(n14753), .ZN(
        n14740) );
  NOR4_X1 U16506 ( .A1(n14742), .A2(n14743), .A3(n14744), .A4(n14745), .ZN(
        n14741) );
  OAI221_X1 U16507 ( .B1(n16381), .B2(n16759), .C1(n16382), .C2(n16753), .A(
        n14755), .ZN(n14752) );
  NAND2_X1 U16508 ( .A1(n14722), .A2(n14723), .ZN(n4947) );
  NOR4_X1 U16509 ( .A1(n14732), .A2(n14733), .A3(n14734), .A4(n14735), .ZN(
        n14722) );
  NOR4_X1 U16510 ( .A1(n14724), .A2(n14725), .A3(n14726), .A4(n14727), .ZN(
        n14723) );
  OAI221_X1 U16511 ( .B1(n16376), .B2(n16759), .C1(n16377), .C2(n16753), .A(
        n14737), .ZN(n14734) );
  NAND2_X1 U16512 ( .A1(n14704), .A2(n14705), .ZN(n4948) );
  NOR4_X1 U16513 ( .A1(n14714), .A2(n14715), .A3(n14716), .A4(n14717), .ZN(
        n14704) );
  NOR4_X1 U16514 ( .A1(n14706), .A2(n14707), .A3(n14708), .A4(n14709), .ZN(
        n14705) );
  OAI221_X1 U16515 ( .B1(n16371), .B2(n16759), .C1(n16372), .C2(n16753), .A(
        n14719), .ZN(n14716) );
  NAND2_X1 U16516 ( .A1(n14686), .A2(n14687), .ZN(n4949) );
  NOR4_X1 U16517 ( .A1(n14696), .A2(n14697), .A3(n14698), .A4(n14699), .ZN(
        n14686) );
  NOR4_X1 U16518 ( .A1(n14688), .A2(n14689), .A3(n14690), .A4(n14691), .ZN(
        n14687) );
  OAI221_X1 U16519 ( .B1(n16366), .B2(n16759), .C1(n16367), .C2(n16753), .A(
        n14701), .ZN(n14698) );
  NAND2_X1 U16520 ( .A1(n14668), .A2(n14669), .ZN(n4950) );
  NOR4_X1 U16521 ( .A1(n14678), .A2(n14679), .A3(n14680), .A4(n14681), .ZN(
        n14668) );
  NOR4_X1 U16522 ( .A1(n14670), .A2(n14671), .A3(n14672), .A4(n14673), .ZN(
        n14669) );
  OAI221_X1 U16523 ( .B1(n16361), .B2(n16759), .C1(n16362), .C2(n16753), .A(
        n14683), .ZN(n14680) );
  NAND2_X1 U16524 ( .A1(n14650), .A2(n14651), .ZN(n4951) );
  NOR4_X1 U16525 ( .A1(n14660), .A2(n14661), .A3(n14662), .A4(n14663), .ZN(
        n14650) );
  NOR4_X1 U16526 ( .A1(n14652), .A2(n14653), .A3(n14654), .A4(n14655), .ZN(
        n14651) );
  OAI221_X1 U16527 ( .B1(n16356), .B2(n16759), .C1(n16357), .C2(n16753), .A(
        n14665), .ZN(n14662) );
  NAND2_X1 U16528 ( .A1(n14632), .A2(n14633), .ZN(n4952) );
  NOR4_X1 U16529 ( .A1(n14642), .A2(n14643), .A3(n14644), .A4(n14645), .ZN(
        n14632) );
  NOR4_X1 U16530 ( .A1(n14634), .A2(n14635), .A3(n14636), .A4(n14637), .ZN(
        n14633) );
  OAI221_X1 U16531 ( .B1(n16351), .B2(n16760), .C1(n16352), .C2(n16754), .A(
        n14647), .ZN(n14644) );
  NAND2_X1 U16532 ( .A1(n14614), .A2(n14615), .ZN(n4953) );
  NOR4_X1 U16533 ( .A1(n14624), .A2(n14625), .A3(n14626), .A4(n14627), .ZN(
        n14614) );
  NOR4_X1 U16534 ( .A1(n14616), .A2(n14617), .A3(n14618), .A4(n14619), .ZN(
        n14615) );
  OAI221_X1 U16535 ( .B1(n16346), .B2(n16760), .C1(n16347), .C2(n16754), .A(
        n14629), .ZN(n14626) );
  NAND2_X1 U16536 ( .A1(n14596), .A2(n14597), .ZN(n4954) );
  NOR4_X1 U16537 ( .A1(n14606), .A2(n14607), .A3(n14608), .A4(n14609), .ZN(
        n14596) );
  NOR4_X1 U16538 ( .A1(n14598), .A2(n14599), .A3(n14600), .A4(n14601), .ZN(
        n14597) );
  OAI221_X1 U16539 ( .B1(n16341), .B2(n16760), .C1(n16342), .C2(n16754), .A(
        n14611), .ZN(n14608) );
  NAND2_X1 U16540 ( .A1(n14578), .A2(n14579), .ZN(n4955) );
  NOR4_X1 U16541 ( .A1(n14588), .A2(n14589), .A3(n14590), .A4(n14591), .ZN(
        n14578) );
  NOR4_X1 U16542 ( .A1(n14580), .A2(n14581), .A3(n14582), .A4(n14583), .ZN(
        n14579) );
  OAI221_X1 U16543 ( .B1(n16336), .B2(n16760), .C1(n16337), .C2(n16754), .A(
        n14593), .ZN(n14590) );
  NAND2_X1 U16544 ( .A1(n14560), .A2(n14561), .ZN(n4956) );
  NOR4_X1 U16545 ( .A1(n14570), .A2(n14571), .A3(n14572), .A4(n14573), .ZN(
        n14560) );
  NOR4_X1 U16546 ( .A1(n14562), .A2(n14563), .A3(n14564), .A4(n14565), .ZN(
        n14561) );
  OAI221_X1 U16547 ( .B1(n16331), .B2(n16760), .C1(n16332), .C2(n16754), .A(
        n14575), .ZN(n14572) );
  NAND2_X1 U16548 ( .A1(n14542), .A2(n14543), .ZN(n4957) );
  NOR4_X1 U16549 ( .A1(n14552), .A2(n14553), .A3(n14554), .A4(n14555), .ZN(
        n14542) );
  NOR4_X1 U16550 ( .A1(n14544), .A2(n14545), .A3(n14546), .A4(n14547), .ZN(
        n14543) );
  OAI221_X1 U16551 ( .B1(n16326), .B2(n16760), .C1(n16327), .C2(n16754), .A(
        n14557), .ZN(n14554) );
  NAND2_X1 U16552 ( .A1(n14524), .A2(n14525), .ZN(n4958) );
  NOR4_X1 U16553 ( .A1(n14534), .A2(n14535), .A3(n14536), .A4(n14537), .ZN(
        n14524) );
  NOR4_X1 U16554 ( .A1(n14526), .A2(n14527), .A3(n14528), .A4(n14529), .ZN(
        n14525) );
  OAI221_X1 U16555 ( .B1(n16321), .B2(n16760), .C1(n16322), .C2(n16754), .A(
        n14539), .ZN(n14536) );
  NAND2_X1 U16556 ( .A1(n14506), .A2(n14507), .ZN(n4959) );
  NOR4_X1 U16557 ( .A1(n14516), .A2(n14517), .A3(n14518), .A4(n14519), .ZN(
        n14506) );
  NOR4_X1 U16558 ( .A1(n14508), .A2(n14509), .A3(n14510), .A4(n14511), .ZN(
        n14507) );
  OAI221_X1 U16559 ( .B1(n16316), .B2(n16760), .C1(n16317), .C2(n16754), .A(
        n14521), .ZN(n14518) );
  NAND2_X1 U16560 ( .A1(n14488), .A2(n14489), .ZN(n4960) );
  NOR4_X1 U16561 ( .A1(n14498), .A2(n14499), .A3(n14500), .A4(n14501), .ZN(
        n14488) );
  NOR4_X1 U16562 ( .A1(n14490), .A2(n14491), .A3(n14492), .A4(n14493), .ZN(
        n14489) );
  OAI221_X1 U16563 ( .B1(n16311), .B2(n16760), .C1(n16312), .C2(n16754), .A(
        n14503), .ZN(n14500) );
  NAND2_X1 U16564 ( .A1(n14470), .A2(n14471), .ZN(n4961) );
  NOR4_X1 U16565 ( .A1(n14480), .A2(n14481), .A3(n14482), .A4(n14483), .ZN(
        n14470) );
  NOR4_X1 U16566 ( .A1(n14472), .A2(n14473), .A3(n14474), .A4(n14475), .ZN(
        n14471) );
  OAI221_X1 U16567 ( .B1(n16306), .B2(n16760), .C1(n16307), .C2(n16754), .A(
        n14485), .ZN(n14482) );
  NAND2_X1 U16568 ( .A1(n14452), .A2(n14453), .ZN(n4962) );
  NOR4_X1 U16569 ( .A1(n14462), .A2(n14463), .A3(n14464), .A4(n14465), .ZN(
        n14452) );
  NOR4_X1 U16570 ( .A1(n14454), .A2(n14455), .A3(n14456), .A4(n14457), .ZN(
        n14453) );
  OAI221_X1 U16571 ( .B1(n16301), .B2(n16760), .C1(n16302), .C2(n16754), .A(
        n14467), .ZN(n14464) );
  NAND2_X1 U16572 ( .A1(n14434), .A2(n14435), .ZN(n4963) );
  NOR4_X1 U16573 ( .A1(n14444), .A2(n14445), .A3(n14446), .A4(n14447), .ZN(
        n14434) );
  NOR4_X1 U16574 ( .A1(n14436), .A2(n14437), .A3(n14438), .A4(n14439), .ZN(
        n14435) );
  OAI221_X1 U16575 ( .B1(n16296), .B2(n16760), .C1(n16297), .C2(n16754), .A(
        n14449), .ZN(n14446) );
  NAND2_X1 U16576 ( .A1(n14416), .A2(n14417), .ZN(n4964) );
  NOR4_X1 U16577 ( .A1(n14426), .A2(n14427), .A3(n14428), .A4(n14429), .ZN(
        n14416) );
  NOR4_X1 U16578 ( .A1(n14418), .A2(n14419), .A3(n14420), .A4(n14421), .ZN(
        n14417) );
  OAI221_X1 U16579 ( .B1(n16291), .B2(n16761), .C1(n16292), .C2(n16755), .A(
        n14431), .ZN(n14428) );
  NAND2_X1 U16580 ( .A1(n14398), .A2(n14399), .ZN(n4965) );
  NOR4_X1 U16581 ( .A1(n14408), .A2(n14409), .A3(n14410), .A4(n14411), .ZN(
        n14398) );
  NOR4_X1 U16582 ( .A1(n14400), .A2(n14401), .A3(n14402), .A4(n14403), .ZN(
        n14399) );
  OAI221_X1 U16583 ( .B1(n16286), .B2(n16761), .C1(n16287), .C2(n16755), .A(
        n14413), .ZN(n14410) );
  NAND2_X1 U16584 ( .A1(n14380), .A2(n14381), .ZN(n4966) );
  NOR4_X1 U16585 ( .A1(n14390), .A2(n14391), .A3(n14392), .A4(n14393), .ZN(
        n14380) );
  NOR4_X1 U16586 ( .A1(n14382), .A2(n14383), .A3(n14384), .A4(n14385), .ZN(
        n14381) );
  OAI221_X1 U16587 ( .B1(n16281), .B2(n16761), .C1(n16282), .C2(n16755), .A(
        n14395), .ZN(n14392) );
  NAND2_X1 U16588 ( .A1(n14362), .A2(n14363), .ZN(n4967) );
  NOR4_X1 U16589 ( .A1(n14372), .A2(n14373), .A3(n14374), .A4(n14375), .ZN(
        n14362) );
  NOR4_X1 U16590 ( .A1(n14364), .A2(n14365), .A3(n14366), .A4(n14367), .ZN(
        n14363) );
  OAI221_X1 U16591 ( .B1(n16276), .B2(n16761), .C1(n16277), .C2(n16755), .A(
        n14377), .ZN(n14374) );
  NAND2_X1 U16592 ( .A1(n14344), .A2(n14345), .ZN(n4968) );
  NOR4_X1 U16593 ( .A1(n14354), .A2(n14355), .A3(n14356), .A4(n14357), .ZN(
        n14344) );
  NOR4_X1 U16594 ( .A1(n14346), .A2(n14347), .A3(n14348), .A4(n14349), .ZN(
        n14345) );
  OAI221_X1 U16595 ( .B1(n16271), .B2(n16761), .C1(n16272), .C2(n16755), .A(
        n14359), .ZN(n14356) );
  NAND2_X1 U16596 ( .A1(n14326), .A2(n14327), .ZN(n4969) );
  NOR4_X1 U16597 ( .A1(n14336), .A2(n14337), .A3(n14338), .A4(n14339), .ZN(
        n14326) );
  NOR4_X1 U16598 ( .A1(n14328), .A2(n14329), .A3(n14330), .A4(n14331), .ZN(
        n14327) );
  OAI221_X1 U16599 ( .B1(n16266), .B2(n16761), .C1(n16267), .C2(n16755), .A(
        n14341), .ZN(n14338) );
  NAND2_X1 U16600 ( .A1(n14308), .A2(n14309), .ZN(n4970) );
  NOR4_X1 U16601 ( .A1(n14318), .A2(n14319), .A3(n14320), .A4(n14321), .ZN(
        n14308) );
  NOR4_X1 U16602 ( .A1(n14310), .A2(n14311), .A3(n14312), .A4(n14313), .ZN(
        n14309) );
  OAI221_X1 U16603 ( .B1(n16261), .B2(n16761), .C1(n16262), .C2(n16755), .A(
        n14323), .ZN(n14320) );
  NAND2_X1 U16604 ( .A1(n14290), .A2(n14291), .ZN(n4971) );
  NOR4_X1 U16605 ( .A1(n14300), .A2(n14301), .A3(n14302), .A4(n14303), .ZN(
        n14290) );
  NOR4_X1 U16606 ( .A1(n14292), .A2(n14293), .A3(n14294), .A4(n14295), .ZN(
        n14291) );
  OAI221_X1 U16607 ( .B1(n16256), .B2(n16761), .C1(n16257), .C2(n16755), .A(
        n14305), .ZN(n14302) );
  NAND2_X1 U16608 ( .A1(n14272), .A2(n14273), .ZN(n4972) );
  NOR4_X1 U16609 ( .A1(n14282), .A2(n14283), .A3(n14284), .A4(n14285), .ZN(
        n14272) );
  NOR4_X1 U16610 ( .A1(n14274), .A2(n14275), .A3(n14276), .A4(n14277), .ZN(
        n14273) );
  OAI221_X1 U16611 ( .B1(n16251), .B2(n16761), .C1(n16252), .C2(n16755), .A(
        n14287), .ZN(n14284) );
  NAND2_X1 U16612 ( .A1(n14254), .A2(n14255), .ZN(n4973) );
  NOR4_X1 U16613 ( .A1(n14264), .A2(n14265), .A3(n14266), .A4(n14267), .ZN(
        n14254) );
  NOR4_X1 U16614 ( .A1(n14256), .A2(n14257), .A3(n14258), .A4(n14259), .ZN(
        n14255) );
  OAI221_X1 U16615 ( .B1(n16246), .B2(n16761), .C1(n16247), .C2(n16755), .A(
        n14269), .ZN(n14266) );
  NAND2_X1 U16616 ( .A1(n14236), .A2(n14237), .ZN(n4974) );
  NOR4_X1 U16617 ( .A1(n14246), .A2(n14247), .A3(n14248), .A4(n14249), .ZN(
        n14236) );
  NOR4_X1 U16618 ( .A1(n14238), .A2(n14239), .A3(n14240), .A4(n14241), .ZN(
        n14237) );
  OAI221_X1 U16619 ( .B1(n16241), .B2(n16761), .C1(n16242), .C2(n16755), .A(
        n14251), .ZN(n14248) );
  NAND2_X1 U16620 ( .A1(n14218), .A2(n14219), .ZN(n4975) );
  NOR4_X1 U16621 ( .A1(n14228), .A2(n14229), .A3(n14230), .A4(n14231), .ZN(
        n14218) );
  NOR4_X1 U16622 ( .A1(n14220), .A2(n14221), .A3(n14222), .A4(n14223), .ZN(
        n14219) );
  OAI221_X1 U16623 ( .B1(n16236), .B2(n16761), .C1(n16237), .C2(n16755), .A(
        n14233), .ZN(n14230) );
  NAND2_X1 U16624 ( .A1(n14200), .A2(n14201), .ZN(n4976) );
  NOR4_X1 U16625 ( .A1(n14210), .A2(n14211), .A3(n14212), .A4(n14213), .ZN(
        n14200) );
  NOR4_X1 U16626 ( .A1(n14202), .A2(n14203), .A3(n14204), .A4(n14205), .ZN(
        n14201) );
  OAI221_X1 U16627 ( .B1(n16231), .B2(n16762), .C1(n16232), .C2(n16756), .A(
        n14215), .ZN(n14212) );
  NAND2_X1 U16628 ( .A1(n14182), .A2(n14183), .ZN(n4977) );
  NOR4_X1 U16629 ( .A1(n14192), .A2(n14193), .A3(n14194), .A4(n14195), .ZN(
        n14182) );
  NOR4_X1 U16630 ( .A1(n14184), .A2(n14185), .A3(n14186), .A4(n14187), .ZN(
        n14183) );
  OAI221_X1 U16631 ( .B1(n16226), .B2(n16762), .C1(n16227), .C2(n16756), .A(
        n14197), .ZN(n14194) );
  NAND2_X1 U16632 ( .A1(n14164), .A2(n14165), .ZN(n4978) );
  NOR4_X1 U16633 ( .A1(n14174), .A2(n14175), .A3(n14176), .A4(n14177), .ZN(
        n14164) );
  NOR4_X1 U16634 ( .A1(n14166), .A2(n14167), .A3(n14168), .A4(n14169), .ZN(
        n14165) );
  OAI221_X1 U16635 ( .B1(n16221), .B2(n16762), .C1(n16222), .C2(n16756), .A(
        n14179), .ZN(n14176) );
  NAND2_X1 U16636 ( .A1(n14146), .A2(n14147), .ZN(n4979) );
  NOR4_X1 U16637 ( .A1(n14156), .A2(n14157), .A3(n14158), .A4(n14159), .ZN(
        n14146) );
  NOR4_X1 U16638 ( .A1(n14148), .A2(n14149), .A3(n14150), .A4(n14151), .ZN(
        n14147) );
  OAI221_X1 U16639 ( .B1(n16216), .B2(n16762), .C1(n16217), .C2(n16756), .A(
        n14161), .ZN(n14158) );
  NAND2_X1 U16640 ( .A1(n14128), .A2(n14129), .ZN(n4980) );
  NOR4_X1 U16641 ( .A1(n14138), .A2(n14139), .A3(n14140), .A4(n14141), .ZN(
        n14128) );
  NOR4_X1 U16642 ( .A1(n14130), .A2(n14131), .A3(n14132), .A4(n14133), .ZN(
        n14129) );
  OAI221_X1 U16643 ( .B1(n16211), .B2(n16762), .C1(n16212), .C2(n16756), .A(
        n14143), .ZN(n14140) );
  NAND2_X1 U16644 ( .A1(n14110), .A2(n14111), .ZN(n4981) );
  NOR4_X1 U16645 ( .A1(n14120), .A2(n14121), .A3(n14122), .A4(n14123), .ZN(
        n14110) );
  NOR4_X1 U16646 ( .A1(n14112), .A2(n14113), .A3(n14114), .A4(n14115), .ZN(
        n14111) );
  OAI221_X1 U16647 ( .B1(n16206), .B2(n16762), .C1(n16207), .C2(n16756), .A(
        n14125), .ZN(n14122) );
  NAND2_X1 U16648 ( .A1(n14092), .A2(n14093), .ZN(n4982) );
  NOR4_X1 U16649 ( .A1(n14102), .A2(n14103), .A3(n14104), .A4(n14105), .ZN(
        n14092) );
  NOR4_X1 U16650 ( .A1(n14094), .A2(n14095), .A3(n14096), .A4(n14097), .ZN(
        n14093) );
  OAI221_X1 U16651 ( .B1(n16201), .B2(n16762), .C1(n16202), .C2(n16756), .A(
        n14107), .ZN(n14104) );
  NAND2_X1 U16652 ( .A1(n14074), .A2(n14075), .ZN(n4983) );
  NOR4_X1 U16653 ( .A1(n14084), .A2(n14085), .A3(n14086), .A4(n14087), .ZN(
        n14074) );
  NOR4_X1 U16654 ( .A1(n14076), .A2(n14077), .A3(n14078), .A4(n14079), .ZN(
        n14075) );
  OAI221_X1 U16655 ( .B1(n16196), .B2(n16762), .C1(n16197), .C2(n16756), .A(
        n14089), .ZN(n14086) );
  NAND2_X1 U16656 ( .A1(n14056), .A2(n14057), .ZN(n4984) );
  NOR4_X1 U16657 ( .A1(n14066), .A2(n14067), .A3(n14068), .A4(n14069), .ZN(
        n14056) );
  NOR4_X1 U16658 ( .A1(n14058), .A2(n14059), .A3(n14060), .A4(n14061), .ZN(
        n14057) );
  OAI221_X1 U16659 ( .B1(n16191), .B2(n16762), .C1(n16192), .C2(n16756), .A(
        n14071), .ZN(n14068) );
  NAND2_X1 U16660 ( .A1(n14038), .A2(n14039), .ZN(n4985) );
  NOR4_X1 U16661 ( .A1(n14048), .A2(n14049), .A3(n14050), .A4(n14051), .ZN(
        n14038) );
  NOR4_X1 U16662 ( .A1(n14040), .A2(n14041), .A3(n14042), .A4(n14043), .ZN(
        n14039) );
  OAI221_X1 U16663 ( .B1(n16186), .B2(n16762), .C1(n16187), .C2(n16756), .A(
        n14053), .ZN(n14050) );
  NAND2_X1 U16664 ( .A1(n14020), .A2(n14021), .ZN(n4986) );
  NOR4_X1 U16665 ( .A1(n14030), .A2(n14031), .A3(n14032), .A4(n14033), .ZN(
        n14020) );
  NOR4_X1 U16666 ( .A1(n14022), .A2(n14023), .A3(n14024), .A4(n14025), .ZN(
        n14021) );
  OAI221_X1 U16667 ( .B1(n16181), .B2(n16762), .C1(n16182), .C2(n16756), .A(
        n14035), .ZN(n14032) );
  NAND2_X1 U16668 ( .A1(n14002), .A2(n14003), .ZN(n4987) );
  NOR4_X1 U16669 ( .A1(n14012), .A2(n14013), .A3(n14014), .A4(n14015), .ZN(
        n14002) );
  NOR4_X1 U16670 ( .A1(n14004), .A2(n14005), .A3(n14006), .A4(n14007), .ZN(
        n14003) );
  OAI221_X1 U16671 ( .B1(n16176), .B2(n16762), .C1(n16177), .C2(n16756), .A(
        n14017), .ZN(n14014) );
  NAND2_X1 U16672 ( .A1(n14976), .A2(n14977), .ZN(n4936) );
  NOR4_X1 U16673 ( .A1(n14986), .A2(n14987), .A3(n14988), .A4(n14989), .ZN(
        n14976) );
  NOR4_X1 U16674 ( .A1(n14978), .A2(n14979), .A3(n14980), .A4(n14981), .ZN(
        n14977) );
  OAI221_X1 U16675 ( .B1(n13446), .B2(n16535), .C1(n968), .C2(n16529), .A(
        n14992), .ZN(n14987) );
  NAND2_X1 U16676 ( .A1(n14958), .A2(n14959), .ZN(n4937) );
  NOR4_X1 U16677 ( .A1(n14968), .A2(n14969), .A3(n14970), .A4(n14971), .ZN(
        n14958) );
  NOR4_X1 U16678 ( .A1(n14960), .A2(n14961), .A3(n14962), .A4(n14963), .ZN(
        n14959) );
  OAI221_X1 U16679 ( .B1(n13445), .B2(n16535), .C1(n967), .C2(n16529), .A(
        n14974), .ZN(n14969) );
  NAND2_X1 U16680 ( .A1(n14940), .A2(n14941), .ZN(n4938) );
  NOR4_X1 U16681 ( .A1(n14950), .A2(n14951), .A3(n14952), .A4(n14953), .ZN(
        n14940) );
  NOR4_X1 U16682 ( .A1(n14942), .A2(n14943), .A3(n14944), .A4(n14945), .ZN(
        n14941) );
  OAI221_X1 U16683 ( .B1(n13444), .B2(n16535), .C1(n966), .C2(n16529), .A(
        n14956), .ZN(n14951) );
  NAND2_X1 U16684 ( .A1(n14888), .A2(n14889), .ZN(n4939) );
  NOR4_X1 U16685 ( .A1(n14915), .A2(n14916), .A3(n14917), .A4(n14918), .ZN(
        n14888) );
  NOR4_X1 U16686 ( .A1(n14890), .A2(n14891), .A3(n14892), .A4(n14893), .ZN(
        n14889) );
  OAI221_X1 U16687 ( .B1(n13443), .B2(n16535), .C1(n965), .C2(n16529), .A(
        n14931), .ZN(n14916) );
  NAND2_X1 U16688 ( .A1(n13768), .A2(n13769), .ZN(n5000) );
  NOR4_X1 U16689 ( .A1(n13778), .A2(n13779), .A3(n13780), .A4(n13781), .ZN(
        n13768) );
  NOR4_X1 U16690 ( .A1(n13770), .A2(n13771), .A3(n13772), .A4(n13773), .ZN(
        n13769) );
  OAI221_X1 U16691 ( .B1(n13446), .B2(n16740), .C1(n968), .C2(n16734), .A(
        n13784), .ZN(n13779) );
  NAND2_X1 U16692 ( .A1(n13750), .A2(n13751), .ZN(n5001) );
  NOR4_X1 U16693 ( .A1(n13760), .A2(n13761), .A3(n13762), .A4(n13763), .ZN(
        n13750) );
  NOR4_X1 U16694 ( .A1(n13752), .A2(n13753), .A3(n13754), .A4(n13755), .ZN(
        n13751) );
  OAI221_X1 U16695 ( .B1(n13445), .B2(n16740), .C1(n967), .C2(n16734), .A(
        n13766), .ZN(n13761) );
  NAND2_X1 U16696 ( .A1(n13732), .A2(n13733), .ZN(n5002) );
  NOR4_X1 U16697 ( .A1(n13742), .A2(n13743), .A3(n13744), .A4(n13745), .ZN(
        n13732) );
  NOR4_X1 U16698 ( .A1(n13734), .A2(n13735), .A3(n13736), .A4(n13737), .ZN(
        n13733) );
  OAI221_X1 U16699 ( .B1(n13444), .B2(n16740), .C1(n966), .C2(n16734), .A(
        n13748), .ZN(n13743) );
  NAND2_X1 U16700 ( .A1(n13680), .A2(n13681), .ZN(n5003) );
  NOR4_X1 U16701 ( .A1(n13707), .A2(n13708), .A3(n13709), .A4(n13710), .ZN(
        n13680) );
  NOR4_X1 U16702 ( .A1(n13682), .A2(n13683), .A3(n13684), .A4(n13685), .ZN(
        n13681) );
  OAI221_X1 U16703 ( .B1(n13443), .B2(n16740), .C1(n965), .C2(n16734), .A(
        n13723), .ZN(n13708) );
  NAND2_X1 U16704 ( .A1(n15192), .A2(n15193), .ZN(n4924) );
  NOR4_X1 U16705 ( .A1(n15202), .A2(n15203), .A3(n15204), .A4(n15205), .ZN(
        n15192) );
  NOR4_X1 U16706 ( .A1(n15194), .A2(n15195), .A3(n15196), .A4(n15197), .ZN(
        n15193) );
  OAI221_X1 U16707 ( .B1(n13458), .B2(n16534), .C1(n980), .C2(n16528), .A(
        n15208), .ZN(n15203) );
  NAND2_X1 U16708 ( .A1(n15174), .A2(n15175), .ZN(n4925) );
  NOR4_X1 U16709 ( .A1(n15184), .A2(n15185), .A3(n15186), .A4(n15187), .ZN(
        n15174) );
  NOR4_X1 U16710 ( .A1(n15176), .A2(n15177), .A3(n15178), .A4(n15179), .ZN(
        n15175) );
  OAI221_X1 U16711 ( .B1(n13457), .B2(n16534), .C1(n979), .C2(n16528), .A(
        n15190), .ZN(n15185) );
  NAND2_X1 U16712 ( .A1(n15156), .A2(n15157), .ZN(n4926) );
  NOR4_X1 U16713 ( .A1(n15166), .A2(n15167), .A3(n15168), .A4(n15169), .ZN(
        n15156) );
  NOR4_X1 U16714 ( .A1(n15158), .A2(n15159), .A3(n15160), .A4(n15161), .ZN(
        n15157) );
  OAI221_X1 U16715 ( .B1(n13456), .B2(n16534), .C1(n978), .C2(n16528), .A(
        n15172), .ZN(n15167) );
  NAND2_X1 U16716 ( .A1(n15138), .A2(n15139), .ZN(n4927) );
  NOR4_X1 U16717 ( .A1(n15148), .A2(n15149), .A3(n15150), .A4(n15151), .ZN(
        n15138) );
  NOR4_X1 U16718 ( .A1(n15140), .A2(n15141), .A3(n15142), .A4(n15143), .ZN(
        n15139) );
  OAI221_X1 U16719 ( .B1(n13455), .B2(n16534), .C1(n977), .C2(n16528), .A(
        n15154), .ZN(n15149) );
  NAND2_X1 U16720 ( .A1(n15120), .A2(n15121), .ZN(n4928) );
  NOR4_X1 U16721 ( .A1(n15130), .A2(n15131), .A3(n15132), .A4(n15133), .ZN(
        n15120) );
  NOR4_X1 U16722 ( .A1(n15122), .A2(n15123), .A3(n15124), .A4(n15125), .ZN(
        n15121) );
  OAI221_X1 U16723 ( .B1(n13454), .B2(n16534), .C1(n976), .C2(n16528), .A(
        n15136), .ZN(n15131) );
  NAND2_X1 U16724 ( .A1(n15102), .A2(n15103), .ZN(n4929) );
  NOR4_X1 U16725 ( .A1(n15112), .A2(n15113), .A3(n15114), .A4(n15115), .ZN(
        n15102) );
  NOR4_X1 U16726 ( .A1(n15104), .A2(n15105), .A3(n15106), .A4(n15107), .ZN(
        n15103) );
  OAI221_X1 U16727 ( .B1(n13453), .B2(n16534), .C1(n975), .C2(n16528), .A(
        n15118), .ZN(n15113) );
  NAND2_X1 U16728 ( .A1(n15084), .A2(n15085), .ZN(n4930) );
  NOR4_X1 U16729 ( .A1(n15094), .A2(n15095), .A3(n15096), .A4(n15097), .ZN(
        n15084) );
  NOR4_X1 U16730 ( .A1(n15086), .A2(n15087), .A3(n15088), .A4(n15089), .ZN(
        n15085) );
  OAI221_X1 U16731 ( .B1(n13452), .B2(n16534), .C1(n974), .C2(n16528), .A(
        n15100), .ZN(n15095) );
  NAND2_X1 U16732 ( .A1(n15066), .A2(n15067), .ZN(n4931) );
  NOR4_X1 U16733 ( .A1(n15076), .A2(n15077), .A3(n15078), .A4(n15079), .ZN(
        n15066) );
  NOR4_X1 U16734 ( .A1(n15068), .A2(n15069), .A3(n15070), .A4(n15071), .ZN(
        n15067) );
  OAI221_X1 U16735 ( .B1(n13451), .B2(n16534), .C1(n973), .C2(n16528), .A(
        n15082), .ZN(n15077) );
  NAND2_X1 U16736 ( .A1(n15048), .A2(n15049), .ZN(n4932) );
  NOR4_X1 U16737 ( .A1(n15058), .A2(n15059), .A3(n15060), .A4(n15061), .ZN(
        n15048) );
  NOR4_X1 U16738 ( .A1(n15050), .A2(n15051), .A3(n15052), .A4(n15053), .ZN(
        n15049) );
  OAI221_X1 U16739 ( .B1(n13450), .B2(n16534), .C1(n972), .C2(n16528), .A(
        n15064), .ZN(n15059) );
  NAND2_X1 U16740 ( .A1(n15030), .A2(n15031), .ZN(n4933) );
  NOR4_X1 U16741 ( .A1(n15040), .A2(n15041), .A3(n15042), .A4(n15043), .ZN(
        n15030) );
  NOR4_X1 U16742 ( .A1(n15032), .A2(n15033), .A3(n15034), .A4(n15035), .ZN(
        n15031) );
  OAI221_X1 U16743 ( .B1(n13449), .B2(n16534), .C1(n971), .C2(n16528), .A(
        n15046), .ZN(n15041) );
  NAND2_X1 U16744 ( .A1(n15012), .A2(n15013), .ZN(n4934) );
  NOR4_X1 U16745 ( .A1(n15022), .A2(n15023), .A3(n15024), .A4(n15025), .ZN(
        n15012) );
  NOR4_X1 U16746 ( .A1(n15014), .A2(n15015), .A3(n15016), .A4(n15017), .ZN(
        n15013) );
  OAI221_X1 U16747 ( .B1(n13448), .B2(n16534), .C1(n970), .C2(n16528), .A(
        n15028), .ZN(n15023) );
  NAND2_X1 U16748 ( .A1(n14994), .A2(n14995), .ZN(n4935) );
  NOR4_X1 U16749 ( .A1(n15004), .A2(n15005), .A3(n15006), .A4(n15007), .ZN(
        n14994) );
  NOR4_X1 U16750 ( .A1(n14996), .A2(n14997), .A3(n14998), .A4(n14999), .ZN(
        n14995) );
  OAI221_X1 U16751 ( .B1(n13447), .B2(n16534), .C1(n969), .C2(n16528), .A(
        n15010), .ZN(n15005) );
  NAND2_X1 U16752 ( .A1(n13984), .A2(n13985), .ZN(n4988) );
  NOR4_X1 U16753 ( .A1(n13994), .A2(n13995), .A3(n13996), .A4(n13997), .ZN(
        n13984) );
  NOR4_X1 U16754 ( .A1(n13986), .A2(n13987), .A3(n13988), .A4(n13989), .ZN(
        n13985) );
  OAI221_X1 U16755 ( .B1(n13458), .B2(n16739), .C1(n980), .C2(n16733), .A(
        n14000), .ZN(n13995) );
  NAND2_X1 U16756 ( .A1(n13966), .A2(n13967), .ZN(n4989) );
  NOR4_X1 U16757 ( .A1(n13976), .A2(n13977), .A3(n13978), .A4(n13979), .ZN(
        n13966) );
  NOR4_X1 U16758 ( .A1(n13968), .A2(n13969), .A3(n13970), .A4(n13971), .ZN(
        n13967) );
  OAI221_X1 U16759 ( .B1(n13457), .B2(n16739), .C1(n979), .C2(n16733), .A(
        n13982), .ZN(n13977) );
  NAND2_X1 U16760 ( .A1(n13948), .A2(n13949), .ZN(n4990) );
  NOR4_X1 U16761 ( .A1(n13958), .A2(n13959), .A3(n13960), .A4(n13961), .ZN(
        n13948) );
  NOR4_X1 U16762 ( .A1(n13950), .A2(n13951), .A3(n13952), .A4(n13953), .ZN(
        n13949) );
  OAI221_X1 U16763 ( .B1(n13456), .B2(n16739), .C1(n978), .C2(n16733), .A(
        n13964), .ZN(n13959) );
  NAND2_X1 U16764 ( .A1(n13930), .A2(n13931), .ZN(n4991) );
  NOR4_X1 U16765 ( .A1(n13940), .A2(n13941), .A3(n13942), .A4(n13943), .ZN(
        n13930) );
  NOR4_X1 U16766 ( .A1(n13932), .A2(n13933), .A3(n13934), .A4(n13935), .ZN(
        n13931) );
  OAI221_X1 U16767 ( .B1(n13455), .B2(n16739), .C1(n977), .C2(n16733), .A(
        n13946), .ZN(n13941) );
  NAND2_X1 U16768 ( .A1(n13912), .A2(n13913), .ZN(n4992) );
  NOR4_X1 U16769 ( .A1(n13922), .A2(n13923), .A3(n13924), .A4(n13925), .ZN(
        n13912) );
  NOR4_X1 U16770 ( .A1(n13914), .A2(n13915), .A3(n13916), .A4(n13917), .ZN(
        n13913) );
  OAI221_X1 U16771 ( .B1(n13454), .B2(n16739), .C1(n976), .C2(n16733), .A(
        n13928), .ZN(n13923) );
  NAND2_X1 U16772 ( .A1(n13894), .A2(n13895), .ZN(n4993) );
  NOR4_X1 U16773 ( .A1(n13904), .A2(n13905), .A3(n13906), .A4(n13907), .ZN(
        n13894) );
  NOR4_X1 U16774 ( .A1(n13896), .A2(n13897), .A3(n13898), .A4(n13899), .ZN(
        n13895) );
  OAI221_X1 U16775 ( .B1(n13453), .B2(n16739), .C1(n975), .C2(n16733), .A(
        n13910), .ZN(n13905) );
  NAND2_X1 U16776 ( .A1(n13876), .A2(n13877), .ZN(n4994) );
  NOR4_X1 U16777 ( .A1(n13886), .A2(n13887), .A3(n13888), .A4(n13889), .ZN(
        n13876) );
  NOR4_X1 U16778 ( .A1(n13878), .A2(n13879), .A3(n13880), .A4(n13881), .ZN(
        n13877) );
  OAI221_X1 U16779 ( .B1(n13452), .B2(n16739), .C1(n974), .C2(n16733), .A(
        n13892), .ZN(n13887) );
  NAND2_X1 U16780 ( .A1(n13858), .A2(n13859), .ZN(n4995) );
  NOR4_X1 U16781 ( .A1(n13868), .A2(n13869), .A3(n13870), .A4(n13871), .ZN(
        n13858) );
  NOR4_X1 U16782 ( .A1(n13860), .A2(n13861), .A3(n13862), .A4(n13863), .ZN(
        n13859) );
  OAI221_X1 U16783 ( .B1(n13451), .B2(n16739), .C1(n973), .C2(n16733), .A(
        n13874), .ZN(n13869) );
  NAND2_X1 U16784 ( .A1(n13840), .A2(n13841), .ZN(n4996) );
  NOR4_X1 U16785 ( .A1(n13850), .A2(n13851), .A3(n13852), .A4(n13853), .ZN(
        n13840) );
  NOR4_X1 U16786 ( .A1(n13842), .A2(n13843), .A3(n13844), .A4(n13845), .ZN(
        n13841) );
  OAI221_X1 U16787 ( .B1(n13450), .B2(n16739), .C1(n972), .C2(n16733), .A(
        n13856), .ZN(n13851) );
  NAND2_X1 U16788 ( .A1(n13822), .A2(n13823), .ZN(n4997) );
  NOR4_X1 U16789 ( .A1(n13832), .A2(n13833), .A3(n13834), .A4(n13835), .ZN(
        n13822) );
  NOR4_X1 U16790 ( .A1(n13824), .A2(n13825), .A3(n13826), .A4(n13827), .ZN(
        n13823) );
  OAI221_X1 U16791 ( .B1(n13449), .B2(n16739), .C1(n971), .C2(n16733), .A(
        n13838), .ZN(n13833) );
  NAND2_X1 U16792 ( .A1(n13804), .A2(n13805), .ZN(n4998) );
  NOR4_X1 U16793 ( .A1(n13814), .A2(n13815), .A3(n13816), .A4(n13817), .ZN(
        n13804) );
  NOR4_X1 U16794 ( .A1(n13806), .A2(n13807), .A3(n13808), .A4(n13809), .ZN(
        n13805) );
  OAI221_X1 U16795 ( .B1(n13448), .B2(n16739), .C1(n970), .C2(n16733), .A(
        n13820), .ZN(n13815) );
  NAND2_X1 U16796 ( .A1(n13786), .A2(n13787), .ZN(n4999) );
  NOR4_X1 U16797 ( .A1(n13796), .A2(n13797), .A3(n13798), .A4(n13799), .ZN(
        n13786) );
  NOR4_X1 U16798 ( .A1(n13788), .A2(n13789), .A3(n13790), .A4(n13791), .ZN(
        n13787) );
  OAI221_X1 U16799 ( .B1(n13447), .B2(n16739), .C1(n969), .C2(n16733), .A(
        n13802), .ZN(n13797) );
  OAI22_X1 U16800 ( .A1(n17234), .A2(n17433), .B1(n17232), .B2(n12709), .ZN(
        n6284) );
  OAI22_X1 U16801 ( .A1(n17234), .A2(n17435), .B1(n17232), .B2(n12708), .ZN(
        n6285) );
  OAI22_X1 U16802 ( .A1(n17234), .A2(n17437), .B1(n17232), .B2(n12707), .ZN(
        n6286) );
  OAI22_X1 U16803 ( .A1(n17234), .A2(n17439), .B1(n17232), .B2(n12706), .ZN(
        n6287) );
  OAI22_X1 U16804 ( .A1(n17234), .A2(n17441), .B1(n17232), .B2(n12705), .ZN(
        n6288) );
  OAI22_X1 U16805 ( .A1(n17235), .A2(n17443), .B1(n17232), .B2(n12704), .ZN(
        n6289) );
  OAI22_X1 U16806 ( .A1(n17235), .A2(n17445), .B1(n17232), .B2(n12703), .ZN(
        n6290) );
  OAI22_X1 U16807 ( .A1(n17235), .A2(n17447), .B1(n17232), .B2(n12702), .ZN(
        n6291) );
  OAI22_X1 U16808 ( .A1(n17235), .A2(n17449), .B1(n17232), .B2(n12701), .ZN(
        n6292) );
  OAI22_X1 U16809 ( .A1(n17235), .A2(n17451), .B1(n17232), .B2(n12700), .ZN(
        n6293) );
  OAI22_X1 U16810 ( .A1(n17236), .A2(n17453), .B1(n17232), .B2(n12699), .ZN(
        n6294) );
  OAI22_X1 U16811 ( .A1(n17236), .A2(n17455), .B1(n17232), .B2(n12698), .ZN(
        n6295) );
  OAI22_X1 U16812 ( .A1(n17236), .A2(n17457), .B1(n17233), .B2(n12697), .ZN(
        n6296) );
  OAI22_X1 U16813 ( .A1(n17236), .A2(n17459), .B1(n17233), .B2(n12696), .ZN(
        n6297) );
  OAI22_X1 U16814 ( .A1(n17236), .A2(n17461), .B1(n17233), .B2(n12695), .ZN(
        n6298) );
  OAI22_X1 U16815 ( .A1(n17237), .A2(n17463), .B1(n17233), .B2(n12694), .ZN(
        n6299) );
  OAI22_X1 U16816 ( .A1(n17237), .A2(n17465), .B1(n17233), .B2(n12693), .ZN(
        n6300) );
  OAI22_X1 U16817 ( .A1(n17237), .A2(n17467), .B1(n17233), .B2(n12692), .ZN(
        n6301) );
  OAI22_X1 U16818 ( .A1(n17237), .A2(n17469), .B1(n17233), .B2(n12691), .ZN(
        n6302) );
  OAI22_X1 U16819 ( .A1(n17237), .A2(n17471), .B1(n17233), .B2(n12690), .ZN(
        n6303) );
  OAI22_X1 U16820 ( .A1(n17238), .A2(n17473), .B1(n17233), .B2(n12689), .ZN(
        n6304) );
  OAI22_X1 U16821 ( .A1(n17238), .A2(n17475), .B1(n17233), .B2(n12688), .ZN(
        n6305) );
  OAI22_X1 U16822 ( .A1(n17238), .A2(n17477), .B1(n17233), .B2(n12687), .ZN(
        n6306) );
  OAI22_X1 U16823 ( .A1(n17238), .A2(n17479), .B1(n17233), .B2(n12686), .ZN(
        n6307) );
  OAI22_X1 U16824 ( .A1(n17238), .A2(n17481), .B1(n17232), .B2(n12685), .ZN(
        n6308) );
  OAI22_X1 U16825 ( .A1(n17239), .A2(n17483), .B1(n17233), .B2(n12684), .ZN(
        n6309) );
  OAI22_X1 U16826 ( .A1(n17239), .A2(n17485), .B1(n17231), .B2(n12683), .ZN(
        n6310) );
  OAI22_X1 U16827 ( .A1(n17239), .A2(n17487), .B1(n17232), .B2(n12682), .ZN(
        n6311) );
  OAI22_X1 U16828 ( .A1(n17239), .A2(n17489), .B1(n17233), .B2(n12681), .ZN(
        n6312) );
  OAI22_X1 U16829 ( .A1(n17239), .A2(n17491), .B1(n17231), .B2(n12680), .ZN(
        n6313) );
  OAI22_X1 U16830 ( .A1(n17240), .A2(n17493), .B1(n17232), .B2(n12679), .ZN(
        n6314) );
  OAI22_X1 U16831 ( .A1(n17240), .A2(n17495), .B1(n17233), .B2(n12678), .ZN(
        n6315) );
  OAI22_X1 U16832 ( .A1(n17240), .A2(n17497), .B1(n17231), .B2(n12677), .ZN(
        n6316) );
  OAI22_X1 U16833 ( .A1(n17240), .A2(n17499), .B1(n17232), .B2(n12676), .ZN(
        n6317) );
  OAI22_X1 U16834 ( .A1(n17240), .A2(n17501), .B1(n17233), .B2(n12675), .ZN(
        n6318) );
  OAI22_X1 U16835 ( .A1(n17241), .A2(n17503), .B1(n17231), .B2(n12674), .ZN(
        n6319) );
  OAI22_X1 U16836 ( .A1(n17241), .A2(n17505), .B1(n13657), .B2(n12673), .ZN(
        n6320) );
  OAI22_X1 U16837 ( .A1(n17241), .A2(n17507), .B1(n17231), .B2(n12672), .ZN(
        n6321) );
  OAI22_X1 U16838 ( .A1(n17241), .A2(n17509), .B1(n13657), .B2(n12671), .ZN(
        n6322) );
  OAI22_X1 U16839 ( .A1(n17241), .A2(n17511), .B1(n17231), .B2(n12670), .ZN(
        n6323) );
  OAI22_X1 U16840 ( .A1(n17242), .A2(n17513), .B1(n13657), .B2(n12669), .ZN(
        n6324) );
  OAI22_X1 U16841 ( .A1(n17242), .A2(n17515), .B1(n17231), .B2(n12668), .ZN(
        n6325) );
  OAI22_X1 U16842 ( .A1(n17242), .A2(n17517), .B1(n17232), .B2(n12667), .ZN(
        n6326) );
  OAI22_X1 U16843 ( .A1(n17242), .A2(n17519), .B1(n17233), .B2(n12666), .ZN(
        n6327) );
  OAI22_X1 U16844 ( .A1(n17242), .A2(n17521), .B1(n17231), .B2(n12665), .ZN(
        n6328) );
  OAI22_X1 U16845 ( .A1(n17243), .A2(n17523), .B1(n17231), .B2(n12664), .ZN(
        n6329) );
  OAI22_X1 U16846 ( .A1(n17243), .A2(n17525), .B1(n17232), .B2(n12663), .ZN(
        n6330) );
  OAI22_X1 U16847 ( .A1(n17243), .A2(n17527), .B1(n17233), .B2(n12662), .ZN(
        n6331) );
  OAI22_X1 U16848 ( .A1(n17243), .A2(n17529), .B1(n17231), .B2(n12661), .ZN(
        n6332) );
  OAI22_X1 U16849 ( .A1(n17243), .A2(n17531), .B1(n17231), .B2(n12660), .ZN(
        n6333) );
  OAI22_X1 U16850 ( .A1(n17244), .A2(n17533), .B1(n13657), .B2(n12659), .ZN(
        n6334) );
  OAI22_X1 U16851 ( .A1(n17244), .A2(n17535), .B1(n17231), .B2(n12658), .ZN(
        n6335) );
  OAI22_X1 U16852 ( .A1(n17244), .A2(n17537), .B1(n13657), .B2(n12657), .ZN(
        n6336) );
  OAI22_X1 U16853 ( .A1(n17244), .A2(n17539), .B1(n17231), .B2(n12656), .ZN(
        n6337) );
  OAI22_X1 U16854 ( .A1(n17244), .A2(n17541), .B1(n13657), .B2(n12655), .ZN(
        n6338) );
  OAI22_X1 U16855 ( .A1(n17245), .A2(n17543), .B1(n17231), .B2(n12654), .ZN(
        n6339) );
  OAI22_X1 U16856 ( .A1(n17245), .A2(n17545), .B1(n13657), .B2(n12653), .ZN(
        n6340) );
  OAI22_X1 U16857 ( .A1(n17245), .A2(n17547), .B1(n17231), .B2(n12652), .ZN(
        n6341) );
  OAI22_X1 U16858 ( .A1(n17245), .A2(n17549), .B1(n13657), .B2(n12651), .ZN(
        n6342) );
  OAI22_X1 U16859 ( .A1(n17245), .A2(n17551), .B1(n17231), .B2(n12650), .ZN(
        n6343) );
  NOR2_X1 U16860 ( .A1(n12196), .A2(ADD_RD2[2]), .ZN(n16065) );
  NOR2_X1 U16861 ( .A1(n12191), .A2(ADD_RD1[2]), .ZN(n14857) );
  NOR2_X1 U16862 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n16066) );
  NOR2_X1 U16863 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n14858) );
  NOR2_X1 U16864 ( .A1(n12195), .A2(ADD_RD2[1]), .ZN(n16073) );
  NOR2_X1 U16865 ( .A1(n12190), .A2(ADD_RD1[1]), .ZN(n14865) );
  NOR3_X1 U16866 ( .A1(n12194), .A2(ADD_RD2[4]), .A3(n12197), .ZN(n16074) );
  NOR3_X1 U16867 ( .A1(n12189), .A2(ADD_RD1[4]), .A3(n12192), .ZN(n14866) );
  NOR3_X1 U16868 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n12194), .ZN(n16068)
         );
  NOR3_X1 U16869 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n12189), .ZN(n14860)
         );
  NOR3_X1 U16870 ( .A1(n12193), .A2(ADD_RD2[3]), .A3(n12197), .ZN(n16067) );
  NOR3_X1 U16871 ( .A1(n12188), .A2(ADD_RD1[3]), .A3(n12192), .ZN(n14859) );
  NOR3_X1 U16872 ( .A1(n12193), .A2(ADD_RD2[0]), .A3(n12194), .ZN(n16063) );
  NOR3_X1 U16873 ( .A1(n12188), .A2(ADD_RD1[0]), .A3(n12189), .ZN(n14855) );
  NOR3_X1 U16874 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n12193), .ZN(n16072)
         );
  NOR3_X1 U16875 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n12188), .ZN(n14864)
         );
  NOR3_X1 U16876 ( .A1(n16560), .A2(RST), .A3(n12180), .ZN(n16064) );
  INV_X1 U16877 ( .A(n16085), .ZN(n12180) );
  NOR3_X1 U16878 ( .A1(n16765), .A2(RST), .A3(n12181), .ZN(n14856) );
  INV_X1 U16879 ( .A(n14877), .ZN(n12181) );
  NAND4_X1 U16880 ( .A1(n16089), .A2(n16090), .A3(n16091), .A4(n16092), .ZN(
        n16085) );
  NOR3_X1 U16881 ( .A1(n16093), .A2(n12182), .A3(n16094), .ZN(n16092) );
  NAND4_X1 U16882 ( .A1(n14881), .A2(n14882), .A3(n14883), .A4(n14884), .ZN(
        n14877) );
  NOR3_X1 U16883 ( .A1(n14885), .A2(n12182), .A3(n14886), .ZN(n14884) );
  INV_X1 U16884 ( .A(ADD_RD2[4]), .ZN(n12193) );
  INV_X1 U16885 ( .A(ADD_RD1[4]), .ZN(n12188) );
  INV_X1 U16886 ( .A(ADD_RD2[3]), .ZN(n12194) );
  INV_X1 U16887 ( .A(ADD_RD1[3]), .ZN(n12189) );
  INV_X1 U16888 ( .A(ADD_RD2[0]), .ZN(n12197) );
  INV_X1 U16889 ( .A(ADD_RD1[0]), .ZN(n12192) );
  AND2_X1 U16890 ( .A1(n17589), .A2(n16095), .ZN(n14923) );
  NAND2_X1 U16891 ( .A1(RD2), .A2(EN), .ZN(n16095) );
  AND2_X1 U16892 ( .A1(n17589), .A2(n14887), .ZN(n13715) );
  NAND2_X1 U16893 ( .A1(RD1), .A2(EN), .ZN(n14887) );
  AND2_X1 U16894 ( .A1(n16087), .A2(ADD_RD2[0]), .ZN(n16083) );
  AND2_X1 U16895 ( .A1(n14879), .A2(ADD_RD1[0]), .ZN(n14875) );
  INV_X1 U16896 ( .A(ADD_RD2[1]), .ZN(n12196) );
  INV_X1 U16897 ( .A(ADD_RD1[1]), .ZN(n12191) );
  AND2_X1 U16898 ( .A1(WR), .A2(EN), .ZN(n13652) );
  INV_X1 U16899 ( .A(ADD_WR[3]), .ZN(n12184) );
  INV_X1 U16900 ( .A(ADD_WR[2]), .ZN(n12185) );
  INV_X1 U16901 ( .A(ADD_WR[0]), .ZN(n12187) );
  INV_X1 U16902 ( .A(ADD_WR[1]), .ZN(n12186) );
  INV_X1 U16903 ( .A(WR), .ZN(n12182) );
  INV_X1 U16904 ( .A(ADD_RD2[2]), .ZN(n12195) );
  INV_X1 U16905 ( .A(ADD_RD1[2]), .ZN(n12190) );
  INV_X1 U16906 ( .A(ADD_WR[4]), .ZN(n12183) );
  INV_X1 U16907 ( .A(RST), .ZN(n12179) );
  CLKBUF_X1 U16908 ( .A(n14939), .Z(n16487) );
  CLKBUF_X1 U16909 ( .A(n14938), .Z(n16493) );
  CLKBUF_X1 U16910 ( .A(n14937), .Z(n16499) );
  CLKBUF_X1 U16911 ( .A(n14935), .Z(n16505) );
  CLKBUF_X1 U16912 ( .A(n14934), .Z(n16511) );
  CLKBUF_X1 U16913 ( .A(n14933), .Z(n16517) );
  CLKBUF_X1 U16914 ( .A(n14932), .Z(n16523) );
  CLKBUF_X1 U16915 ( .A(n14930), .Z(n16529) );
  CLKBUF_X1 U16916 ( .A(n14929), .Z(n16535) );
  CLKBUF_X1 U16917 ( .A(n14928), .Z(n16541) );
  CLKBUF_X1 U16918 ( .A(n14927), .Z(n16547) );
  CLKBUF_X1 U16919 ( .A(n14925), .Z(n16553) );
  CLKBUF_X1 U16920 ( .A(n14924), .Z(n16559) );
  CLKBUF_X1 U16921 ( .A(n14922), .Z(n16570) );
  CLKBUF_X1 U16922 ( .A(n14920), .Z(n16576) );
  CLKBUF_X1 U16923 ( .A(n14919), .Z(n16582) );
  CLKBUF_X1 U16924 ( .A(n14914), .Z(n16588) );
  CLKBUF_X1 U16925 ( .A(n14913), .Z(n16594) );
  CLKBUF_X1 U16926 ( .A(n14912), .Z(n16600) );
  CLKBUF_X1 U16927 ( .A(n14910), .Z(n16606) );
  CLKBUF_X1 U16928 ( .A(n14909), .Z(n16612) );
  CLKBUF_X1 U16929 ( .A(n14908), .Z(n16618) );
  CLKBUF_X1 U16930 ( .A(n14907), .Z(n16624) );
  CLKBUF_X1 U16931 ( .A(n14905), .Z(n16630) );
  CLKBUF_X1 U16932 ( .A(n14904), .Z(n16636) );
  CLKBUF_X1 U16933 ( .A(n14903), .Z(n16642) );
  CLKBUF_X1 U16934 ( .A(n14902), .Z(n16648) );
  CLKBUF_X1 U16935 ( .A(n14900), .Z(n16654) );
  CLKBUF_X1 U16936 ( .A(n14899), .Z(n16660) );
  CLKBUF_X1 U16937 ( .A(n14898), .Z(n16666) );
  CLKBUF_X1 U16938 ( .A(n14897), .Z(n16672) );
  CLKBUF_X1 U16939 ( .A(n14895), .Z(n16678) );
  CLKBUF_X1 U16940 ( .A(n14894), .Z(n16684) );
  CLKBUF_X1 U16941 ( .A(n13731), .Z(n16692) );
  CLKBUF_X1 U16942 ( .A(n13730), .Z(n16698) );
  CLKBUF_X1 U16943 ( .A(n13729), .Z(n16704) );
  CLKBUF_X1 U16944 ( .A(n13727), .Z(n16710) );
  CLKBUF_X1 U16945 ( .A(n13726), .Z(n16716) );
  CLKBUF_X1 U16946 ( .A(n13725), .Z(n16722) );
  CLKBUF_X1 U16947 ( .A(n13724), .Z(n16728) );
  CLKBUF_X1 U16948 ( .A(n13722), .Z(n16734) );
  CLKBUF_X1 U16949 ( .A(n13721), .Z(n16740) );
  CLKBUF_X1 U16950 ( .A(n13720), .Z(n16746) );
  CLKBUF_X1 U16951 ( .A(n13719), .Z(n16752) );
  CLKBUF_X1 U16952 ( .A(n13717), .Z(n16758) );
  CLKBUF_X1 U16953 ( .A(n13716), .Z(n16764) );
  CLKBUF_X1 U16954 ( .A(n13714), .Z(n16775) );
  CLKBUF_X1 U16955 ( .A(n13712), .Z(n16781) );
  CLKBUF_X1 U16956 ( .A(n13711), .Z(n16787) );
  CLKBUF_X1 U16957 ( .A(n13706), .Z(n16793) );
  CLKBUF_X1 U16958 ( .A(n13705), .Z(n16799) );
  CLKBUF_X1 U16959 ( .A(n13704), .Z(n16805) );
  CLKBUF_X1 U16960 ( .A(n13702), .Z(n16811) );
  CLKBUF_X1 U16961 ( .A(n13701), .Z(n16817) );
  CLKBUF_X1 U16962 ( .A(n13700), .Z(n16823) );
  CLKBUF_X1 U16963 ( .A(n13699), .Z(n16829) );
  CLKBUF_X1 U16964 ( .A(n13697), .Z(n16835) );
  CLKBUF_X1 U16965 ( .A(n13696), .Z(n16841) );
  CLKBUF_X1 U16966 ( .A(n13695), .Z(n16847) );
  CLKBUF_X1 U16967 ( .A(n13694), .Z(n16853) );
  CLKBUF_X1 U16968 ( .A(n13692), .Z(n16859) );
  CLKBUF_X1 U16969 ( .A(n13691), .Z(n16865) );
  CLKBUF_X1 U16970 ( .A(n13690), .Z(n16871) );
  CLKBUF_X1 U16971 ( .A(n13689), .Z(n16877) );
  CLKBUF_X1 U16972 ( .A(n13687), .Z(n16883) );
  CLKBUF_X1 U16973 ( .A(n13686), .Z(n16889) );
  CLKBUF_X1 U16974 ( .A(n12179), .Z(n17579) );
  CLKBUF_X1 U16975 ( .A(n12179), .Z(n17580) );
  CLKBUF_X1 U16976 ( .A(n12179), .Z(n17581) );
endmodule

