
module PGNET_NBIT32 ( A, B, Ci, P, G );
  input [31:0] A;
  input [31:0] B;
  output [31:0] P;
  output [31:0] G;
  input Ci;
  wire   Ci;
  assign P[0] = 1'b0;
  assign G[0] = Ci;

  XOR2_X1 U2 ( .A(B[9]), .B(A[9]), .Z(P[9]) );
  XOR2_X1 U3 ( .A(B[8]), .B(A[8]), .Z(P[8]) );
  XOR2_X1 U4 ( .A(B[7]), .B(A[7]), .Z(P[7]) );
  XOR2_X1 U5 ( .A(B[6]), .B(A[6]), .Z(P[6]) );
  XOR2_X1 U6 ( .A(B[5]), .B(A[5]), .Z(P[5]) );
  XOR2_X1 U7 ( .A(B[4]), .B(A[4]), .Z(P[4]) );
  XOR2_X1 U8 ( .A(B[3]), .B(A[3]), .Z(P[3]) );
  XOR2_X1 U9 ( .A(B[31]), .B(A[31]), .Z(P[31]) );
  XOR2_X1 U10 ( .A(B[30]), .B(A[30]), .Z(P[30]) );
  XOR2_X1 U11 ( .A(B[2]), .B(A[2]), .Z(P[2]) );
  XOR2_X1 U12 ( .A(B[29]), .B(A[29]), .Z(P[29]) );
  XOR2_X1 U13 ( .A(B[28]), .B(A[28]), .Z(P[28]) );
  XOR2_X1 U14 ( .A(B[27]), .B(A[27]), .Z(P[27]) );
  XOR2_X1 U15 ( .A(B[26]), .B(A[26]), .Z(P[26]) );
  XOR2_X1 U16 ( .A(B[25]), .B(A[25]), .Z(P[25]) );
  XOR2_X1 U17 ( .A(B[24]), .B(A[24]), .Z(P[24]) );
  XOR2_X1 U18 ( .A(B[23]), .B(A[23]), .Z(P[23]) );
  XOR2_X1 U19 ( .A(B[22]), .B(A[22]), .Z(P[22]) );
  XOR2_X1 U20 ( .A(B[21]), .B(A[21]), .Z(P[21]) );
  XOR2_X1 U21 ( .A(B[20]), .B(A[20]), .Z(P[20]) );
  XOR2_X1 U22 ( .A(B[1]), .B(A[1]), .Z(P[1]) );
  XOR2_X1 U23 ( .A(B[19]), .B(A[19]), .Z(P[19]) );
  XOR2_X1 U24 ( .A(B[18]), .B(A[18]), .Z(P[18]) );
  XOR2_X1 U25 ( .A(B[17]), .B(A[17]), .Z(P[17]) );
  XOR2_X1 U26 ( .A(B[16]), .B(A[16]), .Z(P[16]) );
  XOR2_X1 U27 ( .A(B[15]), .B(A[15]), .Z(P[15]) );
  XOR2_X1 U28 ( .A(B[14]), .B(A[14]), .Z(P[14]) );
  XOR2_X1 U29 ( .A(B[13]), .B(A[13]), .Z(P[13]) );
  XOR2_X1 U30 ( .A(B[12]), .B(A[12]), .Z(P[12]) );
  XOR2_X1 U31 ( .A(B[11]), .B(A[11]), .Z(P[11]) );
  XOR2_X1 U32 ( .A(B[10]), .B(A[10]), .Z(P[10]) );
  AND2_X1 U33 ( .A1(B[9]), .A2(A[9]), .ZN(G[9]) );
  AND2_X1 U34 ( .A1(B[8]), .A2(A[8]), .ZN(G[8]) );
  AND2_X1 U35 ( .A1(B[7]), .A2(A[7]), .ZN(G[7]) );
  AND2_X1 U36 ( .A1(B[6]), .A2(A[6]), .ZN(G[6]) );
  AND2_X1 U37 ( .A1(B[5]), .A2(A[5]), .ZN(G[5]) );
  AND2_X1 U38 ( .A1(B[4]), .A2(A[4]), .ZN(G[4]) );
  AND2_X1 U39 ( .A1(B[3]), .A2(A[3]), .ZN(G[3]) );
  AND2_X1 U40 ( .A1(B[31]), .A2(A[31]), .ZN(G[31]) );
  AND2_X1 U41 ( .A1(B[30]), .A2(A[30]), .ZN(G[30]) );
  AND2_X1 U42 ( .A1(B[2]), .A2(A[2]), .ZN(G[2]) );
  AND2_X1 U43 ( .A1(B[29]), .A2(A[29]), .ZN(G[29]) );
  AND2_X1 U44 ( .A1(B[28]), .A2(A[28]), .ZN(G[28]) );
  AND2_X1 U45 ( .A1(B[27]), .A2(A[27]), .ZN(G[27]) );
  AND2_X1 U46 ( .A1(B[26]), .A2(A[26]), .ZN(G[26]) );
  AND2_X1 U47 ( .A1(B[25]), .A2(A[25]), .ZN(G[25]) );
  AND2_X1 U48 ( .A1(B[24]), .A2(A[24]), .ZN(G[24]) );
  AND2_X1 U49 ( .A1(B[23]), .A2(A[23]), .ZN(G[23]) );
  AND2_X1 U50 ( .A1(B[22]), .A2(A[22]), .ZN(G[22]) );
  AND2_X1 U51 ( .A1(B[21]), .A2(A[21]), .ZN(G[21]) );
  AND2_X1 U52 ( .A1(B[20]), .A2(A[20]), .ZN(G[20]) );
  AND2_X1 U53 ( .A1(B[1]), .A2(A[1]), .ZN(G[1]) );
  AND2_X1 U54 ( .A1(B[19]), .A2(A[19]), .ZN(G[19]) );
  AND2_X1 U55 ( .A1(B[18]), .A2(A[18]), .ZN(G[18]) );
  AND2_X1 U56 ( .A1(B[17]), .A2(A[17]), .ZN(G[17]) );
  AND2_X1 U57 ( .A1(B[16]), .A2(A[16]), .ZN(G[16]) );
  AND2_X1 U58 ( .A1(B[15]), .A2(A[15]), .ZN(G[15]) );
  AND2_X1 U59 ( .A1(B[14]), .A2(A[14]), .ZN(G[14]) );
  AND2_X1 U60 ( .A1(B[13]), .A2(A[13]), .ZN(G[13]) );
  AND2_X1 U61 ( .A1(B[12]), .A2(A[12]), .ZN(G[12]) );
  AND2_X1 U62 ( .A1(B[11]), .A2(A[11]), .ZN(G[11]) );
  AND2_X1 U63 ( .A1(B[10]), .A2(A[10]), .ZN(G[10]) );
endmodule


module SPARSETREE_NBIT32_RADIX4 ( A, B, Ci, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Ci;
  wire   \s_G[4][31] , \s_G[4][27] , \s_G[3][31] , \s_G[3][23] , \s_G[3][15] ,
         \s_G[2][31] , \s_G[2][27] , \s_G[2][23] , \s_G[2][19] , \s_G[2][15] ,
         \s_G[2][11] , \s_G[2][7] , \s_G[1][31] , \s_G[1][29] , \s_G[1][27] ,
         \s_G[1][25] , \s_G[1][23] , \s_G[1][21] , \s_G[1][19] , \s_G[1][17] ,
         \s_G[1][15] , \s_G[1][13] , \s_G[1][11] , \s_G[1][9] , \s_G[1][7] ,
         \s_G[1][5] , \s_G[1][3] , \s_G[1][1] , \s_G[0][31] , \s_G[0][30] ,
         \s_G[0][29] , \s_G[0][28] , \s_G[0][27] , \s_G[0][26] , \s_G[0][25] ,
         \s_G[0][24] , \s_G[0][23] , \s_G[0][22] , \s_G[0][21] , \s_G[0][20] ,
         \s_G[0][19] , \s_G[0][18] , \s_G[0][17] , \s_G[0][16] , \s_G[0][15] ,
         \s_G[0][14] , \s_G[0][13] , \s_G[0][12] , \s_G[0][11] , \s_G[0][10] ,
         \s_G[0][9] , \s_G[0][8] , \s_G[0][7] , \s_G[0][6] , \s_G[0][5] ,
         \s_G[0][4] , \s_G[0][3] , \s_G[0][2] , \s_G[0][1] , \s_G[0][0] ,
         \s_P[4][31] , \s_P[4][27] , \s_P[3][31] , \s_P[3][23] , \s_P[3][15] ,
         \s_P[2][31] , \s_P[2][27] , \s_P[2][23] , \s_P[2][19] , \s_P[2][15] ,
         \s_P[2][11] , \s_P[2][7] , \s_P[1][31] , \s_P[1][29] , \s_P[1][27] ,
         \s_P[1][25] , \s_P[1][23] , \s_P[1][21] , \s_P[1][19] , \s_P[1][17] ,
         \s_P[1][15] , \s_P[1][13] , \s_P[1][11] , \s_P[1][9] , \s_P[1][7] ,
         \s_P[1][5] , \s_P[1][3] , \s_P[0][31] , \s_P[0][30] , \s_P[0][29] ,
         \s_P[0][28] , \s_P[0][27] , \s_P[0][26] , \s_P[0][25] , \s_P[0][24] ,
         \s_P[0][23] , \s_P[0][22] , \s_P[0][21] , \s_P[0][20] , \s_P[0][19] ,
         \s_P[0][18] , \s_P[0][17] , \s_P[0][16] , \s_P[0][15] , \s_P[0][14] ,
         \s_P[0][13] , \s_P[0][12] , \s_P[0][11] , \s_P[0][10] , \s_P[0][9] ,
         \s_P[0][8] , \s_P[0][7] , \s_P[0][6] , \s_P[0][5] , \s_P[0][4] ,
         \s_P[0][3] , \s_P[0][2] , \s_P[0][1] ;
  wire   SYNOPSYS_UNCONNECTED__0;

  PGNET_NBIT32 PGNETWORK ( .A(A), .B(B), .Ci(Ci), .P({\s_P[0][31] , 
        \s_P[0][30] , \s_P[0][29] , \s_P[0][28] , \s_P[0][27] , \s_P[0][26] , 
        \s_P[0][25] , \s_P[0][24] , \s_P[0][23] , \s_P[0][22] , \s_P[0][21] , 
        \s_P[0][20] , \s_P[0][19] , \s_P[0][18] , \s_P[0][17] , \s_P[0][16] , 
        \s_P[0][15] , \s_P[0][14] , \s_P[0][13] , \s_P[0][12] , \s_P[0][11] , 
        \s_P[0][10] , \s_P[0][9] , \s_P[0][8] , \s_P[0][7] , \s_P[0][6] , 
        \s_P[0][5] , \s_P[0][4] , \s_P[0][3] , \s_P[0][2] , \s_P[0][1] , 
        SYNOPSYS_UNCONNECTED__0}), .G({\s_G[0][31] , \s_G[0][30] , 
        \s_G[0][29] , \s_G[0][28] , \s_G[0][27] , \s_G[0][26] , \s_G[0][25] , 
        \s_G[0][24] , \s_G[0][23] , \s_G[0][22] , \s_G[0][21] , \s_G[0][20] , 
        \s_G[0][19] , \s_G[0][18] , \s_G[0][17] , \s_G[0][16] , \s_G[0][15] , 
        \s_G[0][14] , \s_G[0][13] , \s_G[0][12] , \s_G[0][11] , \s_G[0][10] , 
        \s_G[0][9] , \s_G[0][8] , \s_G[0][7] , \s_G[0][6] , \s_G[0][5] , 
        \s_G[0][4] , \s_G[0][3] , \s_G[0][2] , \s_G[0][1] , \s_G[0][0] }) );
  BLOCKG_0 n_G1_1_1 ( .pik(\s_P[0][1] ), .gik(\s_G[0][1] ), .gk_1j(\s_G[0][0] ), .gij(\s_G[1][1] ) );
  BLOCKPG_0 m_PG1_1_3 ( .pik(\s_P[0][3] ), .gik(\s_G[0][3] ), .gk_1j(
        \s_G[0][2] ), .pk_1j(\s_P[0][2] ), .gij(\s_G[1][3] ), .pij(\s_P[1][3] ) );
  BLOCKPG_26 m_PG1_1_5 ( .pik(\s_P[0][5] ), .gik(\s_G[0][5] ), .gk_1j(
        \s_G[0][4] ), .pk_1j(\s_P[0][4] ), .gij(\s_G[1][5] ), .pij(\s_P[1][5] ) );
  BLOCKPG_25 m_PG1_1_7 ( .pik(\s_P[0][7] ), .gik(\s_G[0][7] ), .gk_1j(
        \s_G[0][6] ), .pk_1j(\s_P[0][6] ), .gij(\s_G[1][7] ), .pij(\s_P[1][7] ) );
  BLOCKPG_24 m_PG1_1_9 ( .pik(\s_P[0][9] ), .gik(\s_G[0][9] ), .gk_1j(
        \s_G[0][8] ), .pk_1j(\s_P[0][8] ), .gij(\s_G[1][9] ), .pij(\s_P[1][9] ) );
  BLOCKPG_23 m_PG1_1_11 ( .pik(\s_P[0][11] ), .gik(\s_G[0][11] ), .gk_1j(
        \s_G[0][10] ), .pk_1j(\s_P[0][10] ), .gij(\s_G[1][11] ), .pij(
        \s_P[1][11] ) );
  BLOCKPG_22 m_PG1_1_13 ( .pik(\s_P[0][13] ), .gik(\s_G[0][13] ), .gk_1j(
        \s_G[0][12] ), .pk_1j(\s_P[0][12] ), .gij(\s_G[1][13] ), .pij(
        \s_P[1][13] ) );
  BLOCKPG_21 m_PG1_1_15 ( .pik(\s_P[0][15] ), .gik(\s_G[0][15] ), .gk_1j(
        \s_G[0][14] ), .pk_1j(\s_P[0][14] ), .gij(\s_G[1][15] ), .pij(
        \s_P[1][15] ) );
  BLOCKPG_20 m_PG1_1_17 ( .pik(\s_P[0][17] ), .gik(\s_G[0][17] ), .gk_1j(
        \s_G[0][16] ), .pk_1j(\s_P[0][16] ), .gij(\s_G[1][17] ), .pij(
        \s_P[1][17] ) );
  BLOCKPG_19 m_PG1_1_19 ( .pik(\s_P[0][19] ), .gik(\s_G[0][19] ), .gk_1j(
        \s_G[0][18] ), .pk_1j(\s_P[0][18] ), .gij(\s_G[1][19] ), .pij(
        \s_P[1][19] ) );
  BLOCKPG_18 m_PG1_1_21 ( .pik(\s_P[0][21] ), .gik(\s_G[0][21] ), .gk_1j(
        \s_G[0][20] ), .pk_1j(\s_P[0][20] ), .gij(\s_G[1][21] ), .pij(
        \s_P[1][21] ) );
  BLOCKPG_17 m_PG1_1_23 ( .pik(\s_P[0][23] ), .gik(\s_G[0][23] ), .gk_1j(
        \s_G[0][22] ), .pk_1j(\s_P[0][22] ), .gij(\s_G[1][23] ), .pij(
        \s_P[1][23] ) );
  BLOCKPG_16 m_PG1_1_25 ( .pik(\s_P[0][25] ), .gik(\s_G[0][25] ), .gk_1j(
        \s_G[0][24] ), .pk_1j(\s_P[0][24] ), .gij(\s_G[1][25] ), .pij(
        \s_P[1][25] ) );
  BLOCKPG_15 m_PG1_1_27 ( .pik(\s_P[0][27] ), .gik(\s_G[0][27] ), .gk_1j(
        \s_G[0][26] ), .pk_1j(\s_P[0][26] ), .gij(\s_G[1][27] ), .pij(
        \s_P[1][27] ) );
  BLOCKPG_14 m_PG1_1_29 ( .pik(\s_P[0][29] ), .gik(\s_G[0][29] ), .gk_1j(
        \s_G[0][28] ), .pk_1j(\s_P[0][28] ), .gij(\s_G[1][29] ), .pij(
        \s_P[1][29] ) );
  BLOCKPG_13 m_PG1_1_31 ( .pik(\s_P[0][31] ), .gik(\s_G[0][31] ), .gk_1j(
        \s_G[0][30] ), .pk_1j(\s_P[0][30] ), .gij(\s_G[1][31] ), .pij(
        \s_P[1][31] ) );
  BLOCKG_8 n_G1_2_3 ( .pik(\s_P[1][3] ), .gik(\s_G[1][3] ), .gk_1j(\s_G[1][1] ), .gij(Co[0]) );
  BLOCKPG_12 m_PG1_2_7 ( .pik(\s_P[1][7] ), .gik(\s_G[1][7] ), .gk_1j(
        \s_G[1][5] ), .pk_1j(\s_P[1][5] ), .gij(\s_G[2][7] ), .pij(\s_P[2][7] ) );
  BLOCKPG_11 m_PG1_2_11 ( .pik(\s_P[1][11] ), .gik(\s_G[1][11] ), .gk_1j(
        \s_G[1][9] ), .pk_1j(\s_P[1][9] ), .gij(\s_G[2][11] ), .pij(
        \s_P[2][11] ) );
  BLOCKPG_10 m_PG1_2_15 ( .pik(\s_P[1][15] ), .gik(\s_G[1][15] ), .gk_1j(
        \s_G[1][13] ), .pk_1j(\s_P[1][13] ), .gij(\s_G[2][15] ), .pij(
        \s_P[2][15] ) );
  BLOCKPG_9 m_PG1_2_19 ( .pik(\s_P[1][19] ), .gik(\s_G[1][19] ), .gk_1j(
        \s_G[1][17] ), .pk_1j(\s_P[1][17] ), .gij(\s_G[2][19] ), .pij(
        \s_P[2][19] ) );
  BLOCKPG_8 m_PG1_2_23 ( .pik(\s_P[1][23] ), .gik(\s_G[1][23] ), .gk_1j(
        \s_G[1][21] ), .pk_1j(\s_P[1][21] ), .gij(\s_G[2][23] ), .pij(
        \s_P[2][23] ) );
  BLOCKPG_7 m_PG1_2_27 ( .pik(\s_P[1][27] ), .gik(\s_G[1][27] ), .gk_1j(
        \s_G[1][25] ), .pk_1j(\s_P[1][25] ), .gij(\s_G[2][27] ), .pij(
        \s_P[2][27] ) );
  BLOCKPG_6 m_PG1_2_31 ( .pik(\s_P[1][31] ), .gik(\s_G[1][31] ), .gk_1j(
        \s_G[1][29] ), .pk_1j(\s_P[1][29] ), .gij(\s_G[2][31] ), .pij(
        \s_P[2][31] ) );
  BLOCKG_7 n_G2_3_7 ( .pik(\s_P[2][7] ), .gik(\s_G[2][7] ), .gk_1j(Co[0]), 
        .gij(Co[1]) );
  BLOCKPG_5 m_PG2_3_15 ( .pik(\s_P[2][15] ), .gik(\s_G[2][15] ), .gk_1j(
        \s_G[2][11] ), .pk_1j(\s_P[2][11] ), .gij(\s_G[3][15] ), .pij(
        \s_P[3][15] ) );
  BLOCKPG_4 m_PG2_3_23 ( .pik(\s_P[2][23] ), .gik(\s_G[2][23] ), .gk_1j(
        \s_G[2][19] ), .pk_1j(\s_P[2][19] ), .gij(\s_G[3][23] ), .pij(
        \s_P[3][23] ) );
  BLOCKPG_3 m_PG2_3_31 ( .pik(\s_P[2][31] ), .gik(\s_G[2][31] ), .gk_1j(
        \s_G[2][27] ), .pk_1j(\s_P[2][27] ), .gij(\s_G[3][31] ), .pij(
        \s_P[3][31] ) );
  BLOCKG_6 n_G2_4_11 ( .pik(\s_P[2][11] ), .gik(\s_G[2][11] ), .gk_1j(Co[1]), 
        .gij(Co[2]) );
  BLOCKG_5 n_G2_4_15 ( .pik(\s_P[3][15] ), .gik(\s_G[3][15] ), .gk_1j(Co[1]), 
        .gij(Co[3]) );
  BLOCKPG_2 m_PG2_4_27 ( .pik(\s_P[2][27] ), .gik(\s_G[2][27] ), .gk_1j(
        \s_G[3][23] ), .pk_1j(\s_P[3][23] ), .gij(\s_G[4][27] ), .pij(
        \s_P[4][27] ) );
  BLOCKPG_1 m_PG2_4_31 ( .pik(\s_P[3][31] ), .gik(\s_G[3][31] ), .gk_1j(
        \s_G[3][23] ), .pk_1j(\s_P[3][23] ), .gij(\s_G[4][31] ), .pij(
        \s_P[4][31] ) );
  BLOCKG_4 n_G2_5_19 ( .pik(\s_P[2][19] ), .gik(\s_G[2][19] ), .gk_1j(Co[3]), 
        .gij(Co[4]) );
  BLOCKG_3 n_G2_5_23 ( .pik(\s_P[3][23] ), .gik(\s_G[3][23] ), .gk_1j(Co[3]), 
        .gij(Co[5]) );
  BLOCKG_2 n_G2_5_27 ( .pik(\s_P[4][27] ), .gik(\s_G[4][27] ), .gk_1j(Co[3]), 
        .gij(Co[6]) );
  BLOCKG_1 n_G2_5_31 ( .pik(\s_P[4][31] ), .gik(\s_G[4][31] ), .gk_1j(Co[3]), 
        .gij(Co[7]) );
endmodule


module SUMGEN_NBIT32_RADIX4 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSB_RADIX4_0 GENi_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(S[31:28])
         );
  CSB_RADIX4_7 GENi_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(S[27:24])
         );
  CSB_RADIX4_6 GENi_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(S[23:20])
         );
  CSB_RADIX4_5 GENi_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(S[19:16])
         );
  CSB_RADIX4_4 GENi_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(S[15:12])
         );
  CSB_RADIX4_3 GENi_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  CSB_RADIX4_2 GENi_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSB_RADIX4_1 GENi_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
endmodule


module P4ADDER_NBIT32 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [6:0] carry_ST;

  SPARSETREE_NBIT32_RADIX4 SPARSETREE0 ( .A(A), .B(B), .Ci(Ci), .Co({Co, 
        carry_ST}) );
  SUMGEN_NBIT32_RADIX4 SUMGEN0 ( .A(A), .B(B), .Ci({carry_ST, Ci}), .S(S) );
endmodule

