
module WINDOWED_REGISTER_FILE_NBIT64_M5_N3_F2 ( CLK, RST, EN, RD1, RD2, WR, 
        ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2, CALL, RET, FILL, SPILL, 
        BUSIN, BUSOUT );
  input [3:0] ADD_WR;
  input [3:0] ADD_RD1;
  input [3:0] ADD_RD2;
  input [63:0] DATAIN;
  output [63:0] OUT1;
  output [63:0] OUT2;
  input [63:0] BUSIN;
  output [63:0] BUSOUT;
  input CLK, RST, EN, RD1, RD2, WR, CALL, RET;
  output FILL, SPILL;
  wire   N208, N209, N210, N332, N333, N334, N433, N434, N435, N555, N556,
         N557, N560, N561, N562, N888, N890, N914, N915, N916, N924, N925,
         N926, N927, \U3/U195/Z_0 , \U3/U195/Z_1 , \U3/U195/Z_2 ,
         \U3/U195/Z_3 , \U3/U196/Z_0 , \U3/U196/Z_1 , \U3/U196/Z_2 ,
         \U3/U196/Z_3 , \U3/U196/Z_4 , \U3/U199/Z_0 , \U3/U199/Z_1 ,
         \U3/U199/Z_2 , \U3/U199/Z_3 , \U3/U200/Z_0 , \U3/U200/Z_1 ,
         \U3/U200/Z_2 , \U3/U200/Z_3 , \U3/U200/Z_4 , \U3/U201/Z_0 ,
         \U3/U201/Z_1 , \U3/U201/Z_2 , \U3/U201/Z_3 , \U3/U201/Z_4 ,
         \U3/U202/Z_0 , \U3/U202/Z_1 , \U3/U202/Z_2 , \U3/U202/Z_3 , n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1250, n1258, n1259, n1260, n1261, n1303, n1315, n1316, n1317, n1318,
         n1322, n1327, n1328, n1330, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, \r631/carry[1] , \r631/carry[2] ,
         \r631/carry[3] , \r631/carry[4] , \sub_128_C208/carry[4] ,
         \r646/carry[4] , \r646/carry[3] , \r646/carry[2] , \r642/carry[4] ,
         \r642/carry[3] , \r642/carry[2] , \r638/carry[4] , \r638/carry[3] ,
         \r638/carry[2] , \r507/carry[4] , \r507/carry[3] , \r507/carry[2] ,
         \r473/carry[3] , \r467/carry[4] , \r467/carry[3] , \r467/carry[2] ,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375;
  wire   [4:0] SWP;
  wire   [4:0] CWP;
  assign \U3/U195/Z_3  = ADD_RD2[3];
  assign \U3/U199/Z_3  = ADD_RD1[3];

  DFF_X1 \COUNT_reg[0]  ( .D(n4830), .CK(CLK), .QN(n1330) );
  DFF_X1 \COUNT_reg[1]  ( .D(n4822), .CK(CLK), .Q(n8309), .QN(n5300) );
  DFF_X1 FILLING_reg ( .D(n8375), .CK(CLK), .Q(FILL), .QN(n1327) );
  DFF_X1 \CWP_reg[4]  ( .D(n4821), .CK(CLK), .Q(CWP[4]), .QN(n1303) );
  DFF_X1 \CWP_reg[0]  ( .D(n4820), .CK(CLK), .Q(N888), .QN(n1318) );
  DFF_X1 \CWP_reg[3]  ( .D(n4817), .CK(CLK), .Q(CWP[3]), .QN(n1315) );
  DFF_X1 \CWP_reg[2]  ( .D(n4818), .CK(CLK), .Q(CWP[2]), .QN(n1316) );
  DFF_X1 \CWP_reg[1]  ( .D(n4819), .CK(CLK), .Q(CWP[1]), .QN(n1317) );
  DFF_X1 SPILLING_reg ( .D(n4823), .CK(CLK), .Q(SPILL), .QN(n1322) );
  DFF_X1 \SWP_reg[4]  ( .D(n4828), .CK(CLK), .Q(SWP[4]), .QN(n1250) );
  DFF_X1 \SWP_reg[1]  ( .D(n4826), .CK(CLK), .Q(SWP[1]), .QN(n1260) );
  DFF_X1 \SWP_reg[0]  ( .D(n4827), .CK(CLK), .Q(n5025), .QN(n1261) );
  DFF_X1 \SWP_reg[2]  ( .D(n4825), .CK(CLK), .Q(SWP[2]), .QN(n1259) );
  DFF_X1 \SWP_reg[3]  ( .D(n4824), .CK(CLK), .Q(SWP[3]), .QN(n1258) );
  DFF_X1 \COUNT_reg[2]  ( .D(n4829), .CK(CLK), .QN(n1328) );
  DFF_X1 \REGISTERS_reg[0][63]  ( .D(n3729), .CK(CLK), .Q(n7925), .QN(n4894)
         );
  DFF_X1 \REGISTERS_reg[0][62]  ( .D(n3730), .CK(CLK), .Q(n7926), .QN(n4893)
         );
  DFF_X1 \REGISTERS_reg[0][61]  ( .D(n3731), .CK(CLK), .Q(n7927), .QN(n4892)
         );
  DFF_X1 \REGISTERS_reg[0][60]  ( .D(n3732), .CK(CLK), .Q(n7928), .QN(n4891)
         );
  DFF_X1 \REGISTERS_reg[0][59]  ( .D(n3733), .CK(CLK), .Q(n7929), .QN(n4890)
         );
  DFF_X1 \REGISTERS_reg[0][58]  ( .D(n3734), .CK(CLK), .Q(n7930), .QN(n4889)
         );
  DFF_X1 \REGISTERS_reg[0][57]  ( .D(n3735), .CK(CLK), .Q(n7931), .QN(n4888)
         );
  DFF_X1 \REGISTERS_reg[0][56]  ( .D(n3736), .CK(CLK), .Q(n7932), .QN(n4887)
         );
  DFF_X1 \REGISTERS_reg[0][55]  ( .D(n3737), .CK(CLK), .Q(n7933), .QN(n4886)
         );
  DFF_X1 \REGISTERS_reg[0][54]  ( .D(n3738), .CK(CLK), .Q(n7934), .QN(n4885)
         );
  DFF_X1 \REGISTERS_reg[0][53]  ( .D(n3739), .CK(CLK), .Q(n7935), .QN(n4884)
         );
  DFF_X1 \REGISTERS_reg[0][52]  ( .D(n3740), .CK(CLK), .Q(n7936), .QN(n4883)
         );
  DFF_X1 \REGISTERS_reg[0][51]  ( .D(n3741), .CK(CLK), .Q(n7937), .QN(n4882)
         );
  DFF_X1 \REGISTERS_reg[0][50]  ( .D(n3742), .CK(CLK), .Q(n7938), .QN(n4881)
         );
  DFF_X1 \REGISTERS_reg[0][49]  ( .D(n3743), .CK(CLK), .Q(n7939), .QN(n4880)
         );
  DFF_X1 \REGISTERS_reg[0][48]  ( .D(n3744), .CK(CLK), .Q(n7940), .QN(n4879)
         );
  DFF_X1 \REGISTERS_reg[0][47]  ( .D(n3745), .CK(CLK), .Q(n7941), .QN(n4878)
         );
  DFF_X1 \REGISTERS_reg[0][46]  ( .D(n3746), .CK(CLK), .Q(n7942), .QN(n4877)
         );
  DFF_X1 \REGISTERS_reg[0][45]  ( .D(n3747), .CK(CLK), .Q(n7943), .QN(n4876)
         );
  DFF_X1 \REGISTERS_reg[0][44]  ( .D(n3748), .CK(CLK), .Q(n7944), .QN(n4875)
         );
  DFF_X1 \REGISTERS_reg[0][43]  ( .D(n3749), .CK(CLK), .Q(n7945), .QN(n4874)
         );
  DFF_X1 \REGISTERS_reg[0][42]  ( .D(n3750), .CK(CLK), .Q(n7946), .QN(n4873)
         );
  DFF_X1 \REGISTERS_reg[0][41]  ( .D(n3751), .CK(CLK), .Q(n7947), .QN(n4872)
         );
  DFF_X1 \REGISTERS_reg[0][40]  ( .D(n3752), .CK(CLK), .Q(n7948), .QN(n4871)
         );
  DFF_X1 \REGISTERS_reg[0][39]  ( .D(n3753), .CK(CLK), .Q(n7949), .QN(n4870)
         );
  DFF_X1 \REGISTERS_reg[0][38]  ( .D(n3754), .CK(CLK), .Q(n7950), .QN(n4869)
         );
  DFF_X1 \REGISTERS_reg[0][37]  ( .D(n3755), .CK(CLK), .Q(n7951), .QN(n4868)
         );
  DFF_X1 \REGISTERS_reg[0][36]  ( .D(n3756), .CK(CLK), .Q(n7952), .QN(n4867)
         );
  DFF_X1 \REGISTERS_reg[0][35]  ( .D(n3757), .CK(CLK), .Q(n7953), .QN(n4866)
         );
  DFF_X1 \REGISTERS_reg[0][34]  ( .D(n3758), .CK(CLK), .Q(n7954), .QN(n4865)
         );
  DFF_X1 \REGISTERS_reg[0][33]  ( .D(n3759), .CK(CLK), .Q(n7955), .QN(n4864)
         );
  DFF_X1 \REGISTERS_reg[0][32]  ( .D(n3760), .CK(CLK), .Q(n7956), .QN(n4863)
         );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n3761), .CK(CLK), .Q(n7957), .QN(n4862)
         );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n3762), .CK(CLK), .Q(n7958), .QN(n4861)
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n3763), .CK(CLK), .Q(n7959), .QN(n4860)
         );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n3764), .CK(CLK), .Q(n7960), .QN(n4859)
         );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n3765), .CK(CLK), .Q(n7961), .QN(n4858)
         );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n3766), .CK(CLK), .Q(n7962), .QN(n4857)
         );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n3767), .CK(CLK), .Q(n7963), .QN(n4856)
         );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n3768), .CK(CLK), .Q(n7964), .QN(n4855)
         );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n3769), .CK(CLK), .Q(n7965), .QN(n4854)
         );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n3770), .CK(CLK), .Q(n7966), .QN(n4853)
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n3771), .CK(CLK), .Q(n7967), .QN(n4852)
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n3772), .CK(CLK), .Q(n7968), .QN(n4851)
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n3773), .CK(CLK), .Q(n7969), .QN(n4850)
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n3774), .CK(CLK), .Q(n7970), .QN(n4849)
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n3775), .CK(CLK), .Q(n7971), .QN(n4848)
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n3776), .CK(CLK), .Q(n7972), .QN(n4847)
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n3777), .CK(CLK), .Q(n7973), .QN(n4846)
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n3778), .CK(CLK), .Q(n7974), .QN(n4845)
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n3779), .CK(CLK), .Q(n7975), .QN(n4844)
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n3780), .CK(CLK), .Q(n7976), .QN(n4843)
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n3781), .CK(CLK), .Q(n7977), .QN(n4842)
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n3782), .CK(CLK), .Q(n7978), .QN(n4841)
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n3783), .CK(CLK), .Q(n7979), .QN(n4840) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n3784), .CK(CLK), .Q(n7980), .QN(n4839) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n3785), .CK(CLK), .Q(n7981), .QN(n4838) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n3786), .CK(CLK), .Q(n7982), .QN(n4837) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n3787), .CK(CLK), .Q(n7983), .QN(n4836) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n3788), .CK(CLK), .Q(n7984), .QN(n4835) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n3789), .CK(CLK), .Q(n7985), .QN(n4834) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n3790), .CK(CLK), .Q(n7986), .QN(n4833) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n3791), .CK(CLK), .Q(n7987), .QN(n4832) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n3792), .CK(CLK), .Q(n7988), .QN(n4831) );
  DFF_X1 \REGISTERS_reg[1][63]  ( .D(n3793), .CK(CLK), .Q(n5299) );
  DFF_X1 \REGISTERS_reg[1][62]  ( .D(n3794), .CK(CLK), .Q(n5298) );
  DFF_X1 \REGISTERS_reg[1][61]  ( .D(n3795), .CK(CLK), .Q(n5297) );
  DFF_X1 \REGISTERS_reg[1][60]  ( .D(n3796), .CK(CLK), .Q(n5296) );
  DFF_X1 \REGISTERS_reg[1][59]  ( .D(n3797), .CK(CLK), .Q(n5295) );
  DFF_X1 \REGISTERS_reg[1][58]  ( .D(n3798), .CK(CLK), .Q(n5294) );
  DFF_X1 \REGISTERS_reg[1][57]  ( .D(n3799), .CK(CLK), .Q(n5293) );
  DFF_X1 \REGISTERS_reg[1][56]  ( .D(n3800), .CK(CLK), .Q(n5292) );
  DFF_X1 \REGISTERS_reg[1][55]  ( .D(n3801), .CK(CLK), .Q(n5291) );
  DFF_X1 \REGISTERS_reg[1][54]  ( .D(n3802), .CK(CLK), .Q(n5290) );
  DFF_X1 \REGISTERS_reg[1][53]  ( .D(n3803), .CK(CLK), .Q(n5289) );
  DFF_X1 \REGISTERS_reg[1][52]  ( .D(n3804), .CK(CLK), .Q(n5288) );
  DFF_X1 \REGISTERS_reg[1][51]  ( .D(n3805), .CK(CLK), .Q(n5287) );
  DFF_X1 \REGISTERS_reg[1][50]  ( .D(n3806), .CK(CLK), .Q(n5286) );
  DFF_X1 \REGISTERS_reg[1][49]  ( .D(n3807), .CK(CLK), .Q(n5285) );
  DFF_X1 \REGISTERS_reg[1][48]  ( .D(n3808), .CK(CLK), .Q(n5284) );
  DFF_X1 \REGISTERS_reg[1][47]  ( .D(n3809), .CK(CLK), .Q(n5283) );
  DFF_X1 \REGISTERS_reg[1][46]  ( .D(n3810), .CK(CLK), .Q(n5282) );
  DFF_X1 \REGISTERS_reg[1][45]  ( .D(n3811), .CK(CLK), .Q(n5281) );
  DFF_X1 \REGISTERS_reg[1][44]  ( .D(n3812), .CK(CLK), .Q(n5280) );
  DFF_X1 \REGISTERS_reg[1][43]  ( .D(n3813), .CK(CLK), .Q(n5279) );
  DFF_X1 \REGISTERS_reg[1][42]  ( .D(n3814), .CK(CLK), .Q(n5278) );
  DFF_X1 \REGISTERS_reg[1][41]  ( .D(n3815), .CK(CLK), .Q(n5277) );
  DFF_X1 \REGISTERS_reg[1][40]  ( .D(n3816), .CK(CLK), .Q(n5276) );
  DFF_X1 \REGISTERS_reg[1][39]  ( .D(n3817), .CK(CLK), .Q(n5275) );
  DFF_X1 \REGISTERS_reg[1][38]  ( .D(n3818), .CK(CLK), .Q(n5274) );
  DFF_X1 \REGISTERS_reg[1][37]  ( .D(n3819), .CK(CLK), .Q(n5273) );
  DFF_X1 \REGISTERS_reg[1][36]  ( .D(n3820), .CK(CLK), .Q(n5272) );
  DFF_X1 \REGISTERS_reg[1][35]  ( .D(n3821), .CK(CLK), .Q(n5271) );
  DFF_X1 \REGISTERS_reg[1][34]  ( .D(n3822), .CK(CLK), .Q(n5270) );
  DFF_X1 \REGISTERS_reg[1][33]  ( .D(n3823), .CK(CLK), .Q(n5269) );
  DFF_X1 \REGISTERS_reg[1][32]  ( .D(n3824), .CK(CLK), .Q(n5268) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n3825), .CK(CLK), .Q(n5267) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n3826), .CK(CLK), .Q(n5266) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n3827), .CK(CLK), .Q(n5265) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n3828), .CK(CLK), .Q(n5264) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n3829), .CK(CLK), .Q(n5263) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n3830), .CK(CLK), .Q(n5262) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n3831), .CK(CLK), .Q(n5261) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n3832), .CK(CLK), .Q(n5260) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n3833), .CK(CLK), .Q(n5259) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n3834), .CK(CLK), .Q(n5258) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n3835), .CK(CLK), .Q(n5257) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n3836), .CK(CLK), .Q(n5256) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n3837), .CK(CLK), .Q(n5255) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n3838), .CK(CLK), .Q(n5254) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n3839), .CK(CLK), .Q(n5253) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n3840), .CK(CLK), .Q(n5252) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n3841), .CK(CLK), .Q(n5251) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n3842), .CK(CLK), .Q(n5250) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n3843), .CK(CLK), .Q(n5249) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n3844), .CK(CLK), .Q(n5248) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n3845), .CK(CLK), .Q(n5247) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n3846), .CK(CLK), .Q(n5246) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n3847), .CK(CLK), .Q(n5245) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n3848), .CK(CLK), .Q(n5244) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n3849), .CK(CLK), .Q(n5243) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n3850), .CK(CLK), .Q(n5242) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n3851), .CK(CLK), .Q(n5241) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n3852), .CK(CLK), .Q(n5240) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n3853), .CK(CLK), .Q(n5239) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n3854), .CK(CLK), .Q(n5238) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n3855), .CK(CLK), .Q(n5237) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n3856), .CK(CLK), .Q(n5236) );
  DFF_X1 \REGISTERS_reg[2][63]  ( .D(n3857), .CK(CLK), .Q(n5024) );
  DFF_X1 \REGISTERS_reg[2][62]  ( .D(n3858), .CK(CLK), .Q(n5023) );
  DFF_X1 \REGISTERS_reg[2][61]  ( .D(n3859), .CK(CLK), .Q(n5022) );
  DFF_X1 \REGISTERS_reg[2][60]  ( .D(n3860), .CK(CLK), .Q(n5021) );
  DFF_X1 \REGISTERS_reg[2][59]  ( .D(n3861), .CK(CLK), .Q(n5020) );
  DFF_X1 \REGISTERS_reg[2][58]  ( .D(n3862), .CK(CLK), .Q(n5019) );
  DFF_X1 \REGISTERS_reg[2][57]  ( .D(n3863), .CK(CLK), .Q(n5018) );
  DFF_X1 \REGISTERS_reg[2][56]  ( .D(n3864), .CK(CLK), .Q(n5017) );
  DFF_X1 \REGISTERS_reg[2][55]  ( .D(n3865), .CK(CLK), .Q(n5016) );
  DFF_X1 \REGISTERS_reg[2][54]  ( .D(n3866), .CK(CLK), .Q(n5015) );
  DFF_X1 \REGISTERS_reg[2][53]  ( .D(n3867), .CK(CLK), .Q(n5014) );
  DFF_X1 \REGISTERS_reg[2][52]  ( .D(n3868), .CK(CLK), .Q(n5013) );
  DFF_X1 \REGISTERS_reg[2][51]  ( .D(n3869), .CK(CLK), .Q(n5012) );
  DFF_X1 \REGISTERS_reg[2][50]  ( .D(n3870), .CK(CLK), .Q(n5011) );
  DFF_X1 \REGISTERS_reg[2][49]  ( .D(n3871), .CK(CLK), .Q(n5010) );
  DFF_X1 \REGISTERS_reg[2][48]  ( .D(n3872), .CK(CLK), .Q(n5009) );
  DFF_X1 \REGISTERS_reg[2][47]  ( .D(n3873), .CK(CLK), .Q(n5008) );
  DFF_X1 \REGISTERS_reg[2][46]  ( .D(n3874), .CK(CLK), .Q(n5007) );
  DFF_X1 \REGISTERS_reg[2][45]  ( .D(n3875), .CK(CLK), .Q(n5006) );
  DFF_X1 \REGISTERS_reg[2][44]  ( .D(n3876), .CK(CLK), .Q(n5005) );
  DFF_X1 \REGISTERS_reg[2][43]  ( .D(n3877), .CK(CLK), .Q(n5004) );
  DFF_X1 \REGISTERS_reg[2][42]  ( .D(n3878), .CK(CLK), .Q(n5003) );
  DFF_X1 \REGISTERS_reg[2][41]  ( .D(n3879), .CK(CLK), .Q(n5002) );
  DFF_X1 \REGISTERS_reg[2][40]  ( .D(n3880), .CK(CLK), .Q(n5001) );
  DFF_X1 \REGISTERS_reg[2][39]  ( .D(n3881), .CK(CLK), .Q(n5000) );
  DFF_X1 \REGISTERS_reg[2][38]  ( .D(n3882), .CK(CLK), .Q(n4999) );
  DFF_X1 \REGISTERS_reg[2][37]  ( .D(n3883), .CK(CLK), .Q(n4998) );
  DFF_X1 \REGISTERS_reg[2][36]  ( .D(n3884), .CK(CLK), .Q(n4997) );
  DFF_X1 \REGISTERS_reg[2][35]  ( .D(n3885), .CK(CLK), .Q(n4996) );
  DFF_X1 \REGISTERS_reg[2][34]  ( .D(n3886), .CK(CLK), .Q(n4995) );
  DFF_X1 \REGISTERS_reg[2][33]  ( .D(n3887), .CK(CLK), .Q(n4994) );
  DFF_X1 \REGISTERS_reg[2][32]  ( .D(n3888), .CK(CLK), .Q(n4993) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n3889), .CK(CLK), .Q(n4992) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n3890), .CK(CLK), .Q(n4991) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n3891), .CK(CLK), .Q(n4990) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n3892), .CK(CLK), .Q(n4989) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n3893), .CK(CLK), .Q(n4988) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n3894), .CK(CLK), .Q(n4987) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n3895), .CK(CLK), .Q(n4986) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n3896), .CK(CLK), .Q(n4985) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n3897), .CK(CLK), .Q(n4984) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n3898), .CK(CLK), .Q(n4983) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n3899), .CK(CLK), .Q(n4982) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n3900), .CK(CLK), .Q(n4981) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n3901), .CK(CLK), .Q(n4980) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n3902), .CK(CLK), .Q(n4979) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n3903), .CK(CLK), .Q(n4978) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n3904), .CK(CLK), .Q(n4977) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n3905), .CK(CLK), .Q(n4976) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n3906), .CK(CLK), .Q(n4975) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n3907), .CK(CLK), .Q(n4974) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n3908), .CK(CLK), .Q(n4973) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n3909), .CK(CLK), .Q(n4972) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n3910), .CK(CLK), .Q(n4971) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n3911), .CK(CLK), .Q(n4970) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n3912), .CK(CLK), .Q(n4969) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n3913), .CK(CLK), .Q(n4968) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n3914), .CK(CLK), .Q(n4967) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n3915), .CK(CLK), .Q(n4966) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n3916), .CK(CLK), .Q(n4965) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n3917), .CK(CLK), .Q(n4964) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n3918), .CK(CLK), .Q(n4963) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n3919), .CK(CLK), .Q(n4962) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n3920), .CK(CLK), .Q(n4961) );
  DFF_X1 \REGISTERS_reg[3][63]  ( .D(n3921), .CK(CLK), .Q(n7989), .QN(n5428)
         );
  DFF_X1 \REGISTERS_reg[3][62]  ( .D(n3922), .CK(CLK), .Q(n7990), .QN(n5427)
         );
  DFF_X1 \REGISTERS_reg[3][61]  ( .D(n3923), .CK(CLK), .Q(n7991), .QN(n5426)
         );
  DFF_X1 \REGISTERS_reg[3][60]  ( .D(n3924), .CK(CLK), .Q(n7992), .QN(n5425)
         );
  DFF_X1 \REGISTERS_reg[3][59]  ( .D(n3925), .CK(CLK), .Q(n7993), .QN(n5424)
         );
  DFF_X1 \REGISTERS_reg[3][58]  ( .D(n3926), .CK(CLK), .Q(n7994), .QN(n5423)
         );
  DFF_X1 \REGISTERS_reg[3][57]  ( .D(n3927), .CK(CLK), .Q(n7995), .QN(n5422)
         );
  DFF_X1 \REGISTERS_reg[3][56]  ( .D(n3928), .CK(CLK), .Q(n7996), .QN(n5421)
         );
  DFF_X1 \REGISTERS_reg[3][55]  ( .D(n3929), .CK(CLK), .Q(n7997), .QN(n5420)
         );
  DFF_X1 \REGISTERS_reg[3][54]  ( .D(n3930), .CK(CLK), .Q(n7998), .QN(n5419)
         );
  DFF_X1 \REGISTERS_reg[3][53]  ( .D(n3931), .CK(CLK), .Q(n7999), .QN(n5418)
         );
  DFF_X1 \REGISTERS_reg[3][52]  ( .D(n3932), .CK(CLK), .Q(n8000), .QN(n5417)
         );
  DFF_X1 \REGISTERS_reg[3][51]  ( .D(n3933), .CK(CLK), .Q(n8001), .QN(n5416)
         );
  DFF_X1 \REGISTERS_reg[3][50]  ( .D(n3934), .CK(CLK), .Q(n8002), .QN(n5415)
         );
  DFF_X1 \REGISTERS_reg[3][49]  ( .D(n3935), .CK(CLK), .Q(n8003), .QN(n5414)
         );
  DFF_X1 \REGISTERS_reg[3][48]  ( .D(n3936), .CK(CLK), .Q(n8004), .QN(n5413)
         );
  DFF_X1 \REGISTERS_reg[3][47]  ( .D(n3937), .CK(CLK), .Q(n8005), .QN(n5412)
         );
  DFF_X1 \REGISTERS_reg[3][46]  ( .D(n3938), .CK(CLK), .Q(n8006), .QN(n5411)
         );
  DFF_X1 \REGISTERS_reg[3][45]  ( .D(n3939), .CK(CLK), .Q(n8007), .QN(n5410)
         );
  DFF_X1 \REGISTERS_reg[3][44]  ( .D(n3940), .CK(CLK), .Q(n8008), .QN(n5409)
         );
  DFF_X1 \REGISTERS_reg[3][43]  ( .D(n3941), .CK(CLK), .Q(n8009), .QN(n5408)
         );
  DFF_X1 \REGISTERS_reg[3][42]  ( .D(n3942), .CK(CLK), .Q(n8010), .QN(n5407)
         );
  DFF_X1 \REGISTERS_reg[3][41]  ( .D(n3943), .CK(CLK), .Q(n8011), .QN(n5406)
         );
  DFF_X1 \REGISTERS_reg[3][40]  ( .D(n3944), .CK(CLK), .Q(n8012), .QN(n5405)
         );
  DFF_X1 \REGISTERS_reg[3][39]  ( .D(n3945), .CK(CLK), .Q(n8013), .QN(n5404)
         );
  DFF_X1 \REGISTERS_reg[3][38]  ( .D(n3946), .CK(CLK), .Q(n8014), .QN(n5403)
         );
  DFF_X1 \REGISTERS_reg[3][37]  ( .D(n3947), .CK(CLK), .Q(n8015), .QN(n5402)
         );
  DFF_X1 \REGISTERS_reg[3][36]  ( .D(n3948), .CK(CLK), .Q(n8016), .QN(n5401)
         );
  DFF_X1 \REGISTERS_reg[3][35]  ( .D(n3949), .CK(CLK), .Q(n8017), .QN(n5400)
         );
  DFF_X1 \REGISTERS_reg[3][34]  ( .D(n3950), .CK(CLK), .Q(n8018), .QN(n5399)
         );
  DFF_X1 \REGISTERS_reg[3][33]  ( .D(n3951), .CK(CLK), .Q(n8019), .QN(n5398)
         );
  DFF_X1 \REGISTERS_reg[3][32]  ( .D(n3952), .CK(CLK), .Q(n8020), .QN(n5397)
         );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n3953), .CK(CLK), .Q(n8021), .QN(n5396)
         );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n3954), .CK(CLK), .Q(n8022), .QN(n5395)
         );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n3955), .CK(CLK), .Q(n8023), .QN(n5394)
         );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n3956), .CK(CLK), .Q(n8024), .QN(n5393)
         );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n3957), .CK(CLK), .Q(n8025), .QN(n5392)
         );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n3958), .CK(CLK), .Q(n8026), .QN(n5391)
         );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n3959), .CK(CLK), .Q(n8027), .QN(n5390)
         );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n3960), .CK(CLK), .Q(n8028), .QN(n5389)
         );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n3961), .CK(CLK), .Q(n8029), .QN(n5388)
         );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n3962), .CK(CLK), .Q(n8030), .QN(n5387)
         );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n3963), .CK(CLK), .Q(n8031), .QN(n5386)
         );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n3964), .CK(CLK), .Q(n8032), .QN(n5385)
         );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n3965), .CK(CLK), .Q(n8033), .QN(n5384)
         );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n3966), .CK(CLK), .Q(n8034), .QN(n5383)
         );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n3967), .CK(CLK), .Q(n8035), .QN(n5382)
         );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n3968), .CK(CLK), .Q(n8036), .QN(n5381)
         );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n3969), .CK(CLK), .Q(n8037), .QN(n5380)
         );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n3970), .CK(CLK), .Q(n8038), .QN(n5379)
         );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n3971), .CK(CLK), .Q(n8039), .QN(n5378)
         );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n3972), .CK(CLK), .Q(n8040), .QN(n5377)
         );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n3973), .CK(CLK), .Q(n8041), .QN(n5376)
         );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n3974), .CK(CLK), .Q(n8042), .QN(n5375)
         );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n3975), .CK(CLK), .Q(n8043), .QN(n5374) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n3976), .CK(CLK), .Q(n8044), .QN(n5373) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n3977), .CK(CLK), .Q(n8045), .QN(n5372) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n3978), .CK(CLK), .Q(n8046), .QN(n5371) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n3979), .CK(CLK), .Q(n8047), .QN(n5370) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n3980), .CK(CLK), .Q(n8048), .QN(n5369) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n3981), .CK(CLK), .Q(n8049), .QN(n5368) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n3982), .CK(CLK), .Q(n8050), .QN(n5367) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n3983), .CK(CLK), .Q(n8051), .QN(n5366) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n3984), .CK(CLK), .Q(n8052), .QN(n5365) );
  DFF_X1 \REGISTERS_reg[4][63]  ( .D(n3985), .CK(CLK), .Q(n8053) );
  DFF_X1 \REGISTERS_reg[4][62]  ( .D(n3986), .CK(CLK), .Q(n8054) );
  DFF_X1 \REGISTERS_reg[4][61]  ( .D(n3987), .CK(CLK), .Q(n8055) );
  DFF_X1 \REGISTERS_reg[4][60]  ( .D(n3988), .CK(CLK), .Q(n8056) );
  DFF_X1 \REGISTERS_reg[4][59]  ( .D(n3989), .CK(CLK), .Q(n8057) );
  DFF_X1 \REGISTERS_reg[4][58]  ( .D(n3990), .CK(CLK), .Q(n8058) );
  DFF_X1 \REGISTERS_reg[4][57]  ( .D(n3991), .CK(CLK), .Q(n8059) );
  DFF_X1 \REGISTERS_reg[4][56]  ( .D(n3992), .CK(CLK), .Q(n8060) );
  DFF_X1 \REGISTERS_reg[4][55]  ( .D(n3993), .CK(CLK), .Q(n8061) );
  DFF_X1 \REGISTERS_reg[4][54]  ( .D(n3994), .CK(CLK), .Q(n8062) );
  DFF_X1 \REGISTERS_reg[4][53]  ( .D(n3995), .CK(CLK), .Q(n8063) );
  DFF_X1 \REGISTERS_reg[4][52]  ( .D(n3996), .CK(CLK), .Q(n8064) );
  DFF_X1 \REGISTERS_reg[4][51]  ( .D(n3997), .CK(CLK), .Q(n8065) );
  DFF_X1 \REGISTERS_reg[4][50]  ( .D(n3998), .CK(CLK), .Q(n8066) );
  DFF_X1 \REGISTERS_reg[4][49]  ( .D(n3999), .CK(CLK), .Q(n8067) );
  DFF_X1 \REGISTERS_reg[4][48]  ( .D(n4000), .CK(CLK), .Q(n8068) );
  DFF_X1 \REGISTERS_reg[4][47]  ( .D(n4001), .CK(CLK), .Q(n8069) );
  DFF_X1 \REGISTERS_reg[4][46]  ( .D(n4002), .CK(CLK), .Q(n8070) );
  DFF_X1 \REGISTERS_reg[4][45]  ( .D(n4003), .CK(CLK), .Q(n8071) );
  DFF_X1 \REGISTERS_reg[4][44]  ( .D(n4004), .CK(CLK), .Q(n8072) );
  DFF_X1 \REGISTERS_reg[4][43]  ( .D(n4005), .CK(CLK), .Q(n8073) );
  DFF_X1 \REGISTERS_reg[4][42]  ( .D(n4006), .CK(CLK), .Q(n8074) );
  DFF_X1 \REGISTERS_reg[4][41]  ( .D(n4007), .CK(CLK), .Q(n8075) );
  DFF_X1 \REGISTERS_reg[4][40]  ( .D(n4008), .CK(CLK), .Q(n8076) );
  DFF_X1 \REGISTERS_reg[4][39]  ( .D(n4009), .CK(CLK), .Q(n8077) );
  DFF_X1 \REGISTERS_reg[4][38]  ( .D(n4010), .CK(CLK), .Q(n8078) );
  DFF_X1 \REGISTERS_reg[4][37]  ( .D(n4011), .CK(CLK), .Q(n8079) );
  DFF_X1 \REGISTERS_reg[4][36]  ( .D(n4012), .CK(CLK), .Q(n8080) );
  DFF_X1 \REGISTERS_reg[4][35]  ( .D(n4013), .CK(CLK), .Q(n8081) );
  DFF_X1 \REGISTERS_reg[4][34]  ( .D(n4014), .CK(CLK), .Q(n8082) );
  DFF_X1 \REGISTERS_reg[4][33]  ( .D(n4015), .CK(CLK), .Q(n8083) );
  DFF_X1 \REGISTERS_reg[4][32]  ( .D(n4016), .CK(CLK), .Q(n8084) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n4017), .CK(CLK), .Q(n8085) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n4018), .CK(CLK), .Q(n8086) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n4019), .CK(CLK), .Q(n8087) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n4020), .CK(CLK), .Q(n8088) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n4021), .CK(CLK), .Q(n8089) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n4022), .CK(CLK), .Q(n8090) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n4023), .CK(CLK), .Q(n8091) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n4024), .CK(CLK), .Q(n8092) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n4025), .CK(CLK), .Q(n8093) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n4026), .CK(CLK), .Q(n8094) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n4027), .CK(CLK), .Q(n8095) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n4028), .CK(CLK), .Q(n8096) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n4029), .CK(CLK), .Q(n8097) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n4030), .CK(CLK), .Q(n8098) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n4031), .CK(CLK), .Q(n8099) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n4032), .CK(CLK), .Q(n8100) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n4033), .CK(CLK), .Q(n8101) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n4034), .CK(CLK), .Q(n8102) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n4035), .CK(CLK), .Q(n8103) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n4036), .CK(CLK), .Q(n8104) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n4037), .CK(CLK), .Q(n8105) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n4038), .CK(CLK), .Q(n8106) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n4039), .CK(CLK), .Q(n8107) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n4040), .CK(CLK), .Q(n8108) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n4041), .CK(CLK), .Q(n8109) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n4042), .CK(CLK), .Q(n8110) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n4043), .CK(CLK), .Q(n8111) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n4044), .CK(CLK), .Q(n8112) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n4045), .CK(CLK), .Q(n8113) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n4046), .CK(CLK), .Q(n8114) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n4047), .CK(CLK), .Q(n8115) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n4048), .CK(CLK), .Q(n8116) );
  DFF_X1 \REGISTERS_reg[5][63]  ( .D(n4049), .CK(CLK), .Q(n5622), .QN(n482) );
  DFF_X1 \REGISTERS_reg[5][62]  ( .D(n4050), .CK(CLK), .Q(n5621), .QN(n483) );
  DFF_X1 \REGISTERS_reg[5][61]  ( .D(n4051), .CK(CLK), .Q(n5620), .QN(n484) );
  DFF_X1 \REGISTERS_reg[5][60]  ( .D(n4052), .CK(CLK), .Q(n5619), .QN(n485) );
  DFF_X1 \REGISTERS_reg[5][59]  ( .D(n4053), .CK(CLK), .Q(n5618), .QN(n486) );
  DFF_X1 \REGISTERS_reg[5][58]  ( .D(n4054), .CK(CLK), .Q(n5617), .QN(n487) );
  DFF_X1 \REGISTERS_reg[5][57]  ( .D(n4055), .CK(CLK), .Q(n5616), .QN(n488) );
  DFF_X1 \REGISTERS_reg[5][56]  ( .D(n4056), .CK(CLK), .Q(n5615), .QN(n489) );
  DFF_X1 \REGISTERS_reg[5][55]  ( .D(n4057), .CK(CLK), .Q(n5614), .QN(n490) );
  DFF_X1 \REGISTERS_reg[5][54]  ( .D(n4058), .CK(CLK), .Q(n5613), .QN(n491) );
  DFF_X1 \REGISTERS_reg[5][53]  ( .D(n4059), .CK(CLK), .Q(n5612), .QN(n492) );
  DFF_X1 \REGISTERS_reg[5][52]  ( .D(n4060), .CK(CLK), .Q(n5611), .QN(n493) );
  DFF_X1 \REGISTERS_reg[5][51]  ( .D(n4061), .CK(CLK), .Q(n5610), .QN(n494) );
  DFF_X1 \REGISTERS_reg[5][50]  ( .D(n4062), .CK(CLK), .Q(n5609), .QN(n495) );
  DFF_X1 \REGISTERS_reg[5][49]  ( .D(n4063), .CK(CLK), .Q(n5608), .QN(n496) );
  DFF_X1 \REGISTERS_reg[5][48]  ( .D(n4064), .CK(CLK), .Q(n5607), .QN(n497) );
  DFF_X1 \REGISTERS_reg[5][47]  ( .D(n4065), .CK(CLK), .Q(n5606), .QN(n498) );
  DFF_X1 \REGISTERS_reg[5][46]  ( .D(n4066), .CK(CLK), .Q(n5605), .QN(n499) );
  DFF_X1 \REGISTERS_reg[5][45]  ( .D(n4067), .CK(CLK), .Q(n5604), .QN(n500) );
  DFF_X1 \REGISTERS_reg[5][44]  ( .D(n4068), .CK(CLK), .Q(n5603), .QN(n501) );
  DFF_X1 \REGISTERS_reg[5][43]  ( .D(n4069), .CK(CLK), .Q(n5602), .QN(n502) );
  DFF_X1 \REGISTERS_reg[5][42]  ( .D(n4070), .CK(CLK), .Q(n5601), .QN(n503) );
  DFF_X1 \REGISTERS_reg[5][41]  ( .D(n4071), .CK(CLK), .Q(n5600), .QN(n504) );
  DFF_X1 \REGISTERS_reg[5][40]  ( .D(n4072), .CK(CLK), .Q(n5599), .QN(n505) );
  DFF_X1 \REGISTERS_reg[5][39]  ( .D(n4073), .CK(CLK), .Q(n5598), .QN(n506) );
  DFF_X1 \REGISTERS_reg[5][38]  ( .D(n4074), .CK(CLK), .Q(n5597), .QN(n507) );
  DFF_X1 \REGISTERS_reg[5][37]  ( .D(n4075), .CK(CLK), .Q(n5596), .QN(n508) );
  DFF_X1 \REGISTERS_reg[5][36]  ( .D(n4076), .CK(CLK), .Q(n5595), .QN(n509) );
  DFF_X1 \REGISTERS_reg[5][35]  ( .D(n4077), .CK(CLK), .Q(n5594), .QN(n510) );
  DFF_X1 \REGISTERS_reg[5][34]  ( .D(n4078), .CK(CLK), .Q(n5593), .QN(n511) );
  DFF_X1 \REGISTERS_reg[5][33]  ( .D(n4079), .CK(CLK), .Q(n5592), .QN(n512) );
  DFF_X1 \REGISTERS_reg[5][32]  ( .D(n4080), .CK(CLK), .Q(n5591), .QN(n513) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n4081), .CK(CLK), .Q(n5590), .QN(n514) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n4082), .CK(CLK), .Q(n5589), .QN(n515) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n4083), .CK(CLK), .Q(n5588), .QN(n516) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n4084), .CK(CLK), .Q(n5587), .QN(n517) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n4085), .CK(CLK), .Q(n5586), .QN(n518) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n4086), .CK(CLK), .Q(n5585), .QN(n519) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n4087), .CK(CLK), .Q(n5584), .QN(n520) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n4088), .CK(CLK), .Q(n5583), .QN(n521) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n4089), .CK(CLK), .Q(n5582), .QN(n522) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n4090), .CK(CLK), .Q(n5581), .QN(n523) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n4091), .CK(CLK), .Q(n5580), .QN(n524) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n4092), .CK(CLK), .Q(n5579), .QN(n525) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n4093), .CK(CLK), .Q(n5578), .QN(n526) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n4094), .CK(CLK), .Q(n5577), .QN(n527) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n4095), .CK(CLK), .Q(n5576), .QN(n528) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n4096), .CK(CLK), .Q(n5575), .QN(n529) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n4097), .CK(CLK), .Q(n5574), .QN(n530) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n4098), .CK(CLK), .Q(n5573), .QN(n531) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n4099), .CK(CLK), .Q(n5572), .QN(n532) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n4100), .CK(CLK), .Q(n5571), .QN(n533) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n4101), .CK(CLK), .Q(n5570), .QN(n534) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n4102), .CK(CLK), .Q(n5569), .QN(n535) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n4103), .CK(CLK), .Q(n5568), .QN(n536) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n4104), .CK(CLK), .Q(n5567), .QN(n537) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n4105), .CK(CLK), .Q(n5566), .QN(n538) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n4106), .CK(CLK), .Q(n5565), .QN(n539) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n4107), .CK(CLK), .Q(n5564), .QN(n540) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n4108), .CK(CLK), .Q(n5563), .QN(n541) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n4109), .CK(CLK), .Q(n5562), .QN(n542) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n4110), .CK(CLK), .Q(n5561), .QN(n543) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n4111), .CK(CLK), .Q(n5560), .QN(n544) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n4112), .CK(CLK), .Q(n5559), .QN(n545) );
  DFF_X1 \REGISTERS_reg[6][63]  ( .D(n4113), .CK(CLK), .Q(n5814), .QN(n546) );
  DFF_X1 \REGISTERS_reg[6][62]  ( .D(n4114), .CK(CLK), .Q(n5813), .QN(n547) );
  DFF_X1 \REGISTERS_reg[6][61]  ( .D(n4115), .CK(CLK), .Q(n5812), .QN(n548) );
  DFF_X1 \REGISTERS_reg[6][60]  ( .D(n4116), .CK(CLK), .Q(n5811), .QN(n549) );
  DFF_X1 \REGISTERS_reg[6][59]  ( .D(n4117), .CK(CLK), .Q(n5810), .QN(n550) );
  DFF_X1 \REGISTERS_reg[6][58]  ( .D(n4118), .CK(CLK), .Q(n5809), .QN(n551) );
  DFF_X1 \REGISTERS_reg[6][57]  ( .D(n4119), .CK(CLK), .Q(n5808), .QN(n552) );
  DFF_X1 \REGISTERS_reg[6][56]  ( .D(n4120), .CK(CLK), .Q(n5807), .QN(n553) );
  DFF_X1 \REGISTERS_reg[6][55]  ( .D(n4121), .CK(CLK), .Q(n5806), .QN(n554) );
  DFF_X1 \REGISTERS_reg[6][54]  ( .D(n4122), .CK(CLK), .Q(n5805), .QN(n555) );
  DFF_X1 \REGISTERS_reg[6][53]  ( .D(n4123), .CK(CLK), .Q(n5804), .QN(n556) );
  DFF_X1 \REGISTERS_reg[6][52]  ( .D(n4124), .CK(CLK), .Q(n5803), .QN(n557) );
  DFF_X1 \REGISTERS_reg[6][51]  ( .D(n4125), .CK(CLK), .Q(n5802), .QN(n558) );
  DFF_X1 \REGISTERS_reg[6][50]  ( .D(n4126), .CK(CLK), .Q(n5801), .QN(n559) );
  DFF_X1 \REGISTERS_reg[6][49]  ( .D(n4127), .CK(CLK), .Q(n5800), .QN(n560) );
  DFF_X1 \REGISTERS_reg[6][48]  ( .D(n4128), .CK(CLK), .Q(n5799), .QN(n561) );
  DFF_X1 \REGISTERS_reg[6][47]  ( .D(n4129), .CK(CLK), .Q(n5798), .QN(n562) );
  DFF_X1 \REGISTERS_reg[6][46]  ( .D(n4130), .CK(CLK), .Q(n5797), .QN(n563) );
  DFF_X1 \REGISTERS_reg[6][45]  ( .D(n4131), .CK(CLK), .Q(n5796), .QN(n564) );
  DFF_X1 \REGISTERS_reg[6][44]  ( .D(n4132), .CK(CLK), .Q(n5795), .QN(n565) );
  DFF_X1 \REGISTERS_reg[6][43]  ( .D(n4133), .CK(CLK), .Q(n5794), .QN(n566) );
  DFF_X1 \REGISTERS_reg[6][42]  ( .D(n4134), .CK(CLK), .Q(n5793), .QN(n567) );
  DFF_X1 \REGISTERS_reg[6][41]  ( .D(n4135), .CK(CLK), .Q(n5792), .QN(n568) );
  DFF_X1 \REGISTERS_reg[6][40]  ( .D(n4136), .CK(CLK), .Q(n5791), .QN(n569) );
  DFF_X1 \REGISTERS_reg[6][39]  ( .D(n4137), .CK(CLK), .Q(n5790), .QN(n570) );
  DFF_X1 \REGISTERS_reg[6][38]  ( .D(n4138), .CK(CLK), .Q(n5789), .QN(n571) );
  DFF_X1 \REGISTERS_reg[6][37]  ( .D(n4139), .CK(CLK), .Q(n5788), .QN(n572) );
  DFF_X1 \REGISTERS_reg[6][36]  ( .D(n4140), .CK(CLK), .Q(n5787), .QN(n573) );
  DFF_X1 \REGISTERS_reg[6][35]  ( .D(n4141), .CK(CLK), .Q(n5786), .QN(n574) );
  DFF_X1 \REGISTERS_reg[6][34]  ( .D(n4142), .CK(CLK), .Q(n5785), .QN(n575) );
  DFF_X1 \REGISTERS_reg[6][33]  ( .D(n4143), .CK(CLK), .Q(n5784), .QN(n576) );
  DFF_X1 \REGISTERS_reg[6][32]  ( .D(n4144), .CK(CLK), .Q(n5783), .QN(n577) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n4145), .CK(CLK), .Q(n5782), .QN(n578) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n4146), .CK(CLK), .Q(n5781), .QN(n579) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n4147), .CK(CLK), .Q(n5780), .QN(n580) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n4148), .CK(CLK), .Q(n5779), .QN(n581) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n4149), .CK(CLK), .Q(n5778), .QN(n582) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n4150), .CK(CLK), .Q(n5777), .QN(n583) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n4151), .CK(CLK), .Q(n5776), .QN(n584) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n4152), .CK(CLK), .Q(n5775), .QN(n585) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n4153), .CK(CLK), .Q(n5774), .QN(n586) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n4154), .CK(CLK), .Q(n5773), .QN(n587) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n4155), .CK(CLK), .Q(n5772), .QN(n588) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n4156), .CK(CLK), .Q(n5771), .QN(n589) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n4157), .CK(CLK), .Q(n5770), .QN(n590) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n4158), .CK(CLK), .Q(n5769), .QN(n591) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n4159), .CK(CLK), .Q(n5768), .QN(n592) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n4160), .CK(CLK), .Q(n5767), .QN(n593) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n4161), .CK(CLK), .Q(n5766), .QN(n594) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n4162), .CK(CLK), .Q(n5765), .QN(n595) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n4163), .CK(CLK), .Q(n5764), .QN(n596) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n4164), .CK(CLK), .Q(n5763), .QN(n597) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n4165), .CK(CLK), .Q(n5762), .QN(n598) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n4166), .CK(CLK), .Q(n5761), .QN(n599) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n4167), .CK(CLK), .Q(n5760), .QN(n600) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n4168), .CK(CLK), .Q(n5759), .QN(n601) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n4169), .CK(CLK), .Q(n5758), .QN(n602) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n4170), .CK(CLK), .Q(n5757), .QN(n603) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n4171), .CK(CLK), .Q(n5756), .QN(n604) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n4172), .CK(CLK), .Q(n5755), .QN(n605) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n4173), .CK(CLK), .Q(n5754), .QN(n606) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n4174), .CK(CLK), .Q(n5753), .QN(n607) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n4175), .CK(CLK), .Q(n5752), .QN(n608) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n4176), .CK(CLK), .Q(n5751), .QN(n609) );
  DFF_X1 \REGISTERS_reg[7][63]  ( .D(n4177), .CK(CLK), .Q(n8117) );
  DFF_X1 \REGISTERS_reg[7][62]  ( .D(n4178), .CK(CLK), .Q(n8118) );
  DFF_X1 \REGISTERS_reg[7][61]  ( .D(n4179), .CK(CLK), .Q(n8119) );
  DFF_X1 \REGISTERS_reg[7][60]  ( .D(n4180), .CK(CLK), .Q(n8120) );
  DFF_X1 \REGISTERS_reg[7][59]  ( .D(n4181), .CK(CLK), .Q(n8121) );
  DFF_X1 \REGISTERS_reg[7][58]  ( .D(n4182), .CK(CLK), .Q(n8122) );
  DFF_X1 \REGISTERS_reg[7][57]  ( .D(n4183), .CK(CLK), .Q(n8123) );
  DFF_X1 \REGISTERS_reg[7][56]  ( .D(n4184), .CK(CLK), .Q(n8124) );
  DFF_X1 \REGISTERS_reg[7][55]  ( .D(n4185), .CK(CLK), .Q(n8125) );
  DFF_X1 \REGISTERS_reg[7][54]  ( .D(n4186), .CK(CLK), .Q(n8126) );
  DFF_X1 \REGISTERS_reg[7][53]  ( .D(n4187), .CK(CLK), .Q(n8127) );
  DFF_X1 \REGISTERS_reg[7][52]  ( .D(n4188), .CK(CLK), .Q(n8128) );
  DFF_X1 \REGISTERS_reg[7][51]  ( .D(n4189), .CK(CLK), .Q(n8129) );
  DFF_X1 \REGISTERS_reg[7][50]  ( .D(n4190), .CK(CLK), .Q(n8130) );
  DFF_X1 \REGISTERS_reg[7][49]  ( .D(n4191), .CK(CLK), .Q(n8131) );
  DFF_X1 \REGISTERS_reg[7][48]  ( .D(n4192), .CK(CLK), .Q(n8132) );
  DFF_X1 \REGISTERS_reg[7][47]  ( .D(n4193), .CK(CLK), .Q(n8133) );
  DFF_X1 \REGISTERS_reg[7][46]  ( .D(n4194), .CK(CLK), .Q(n8134) );
  DFF_X1 \REGISTERS_reg[7][45]  ( .D(n4195), .CK(CLK), .Q(n8135) );
  DFF_X1 \REGISTERS_reg[7][44]  ( .D(n4196), .CK(CLK), .Q(n8136) );
  DFF_X1 \REGISTERS_reg[7][43]  ( .D(n4197), .CK(CLK), .Q(n8137) );
  DFF_X1 \REGISTERS_reg[7][42]  ( .D(n4198), .CK(CLK), .Q(n8138) );
  DFF_X1 \REGISTERS_reg[7][41]  ( .D(n4199), .CK(CLK), .Q(n8139) );
  DFF_X1 \REGISTERS_reg[7][40]  ( .D(n4200), .CK(CLK), .Q(n8140) );
  DFF_X1 \REGISTERS_reg[7][39]  ( .D(n4201), .CK(CLK), .Q(n8141) );
  DFF_X1 \REGISTERS_reg[7][38]  ( .D(n4202), .CK(CLK), .Q(n8142) );
  DFF_X1 \REGISTERS_reg[7][37]  ( .D(n4203), .CK(CLK), .Q(n8143) );
  DFF_X1 \REGISTERS_reg[7][36]  ( .D(n4204), .CK(CLK), .Q(n8144) );
  DFF_X1 \REGISTERS_reg[7][35]  ( .D(n4205), .CK(CLK), .Q(n8145) );
  DFF_X1 \REGISTERS_reg[7][34]  ( .D(n4206), .CK(CLK), .Q(n8146) );
  DFF_X1 \REGISTERS_reg[7][33]  ( .D(n4207), .CK(CLK), .Q(n8147) );
  DFF_X1 \REGISTERS_reg[7][32]  ( .D(n4208), .CK(CLK), .Q(n8148) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n4209), .CK(CLK), .Q(n8149) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n4210), .CK(CLK), .Q(n8150) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n4211), .CK(CLK), .Q(n8151) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n4212), .CK(CLK), .Q(n8152) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n4213), .CK(CLK), .Q(n8153) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n4214), .CK(CLK), .Q(n8154) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n4215), .CK(CLK), .Q(n8155) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n4216), .CK(CLK), .Q(n8156) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n4217), .CK(CLK), .Q(n8157) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n4218), .CK(CLK), .Q(n8158) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n4219), .CK(CLK), .Q(n8159) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n4220), .CK(CLK), .Q(n8160) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n4221), .CK(CLK), .Q(n8161) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n4222), .CK(CLK), .Q(n8162) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n4223), .CK(CLK), .Q(n8163) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n4224), .CK(CLK), .Q(n8164) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n4225), .CK(CLK), .Q(n8165) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n4226), .CK(CLK), .Q(n8166) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n4227), .CK(CLK), .Q(n8167) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n4228), .CK(CLK), .Q(n8168) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n4229), .CK(CLK), .Q(n8169) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n4230), .CK(CLK), .Q(n8170) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n4231), .CK(CLK), .Q(n8171) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n4232), .CK(CLK), .Q(n8172) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n4233), .CK(CLK), .Q(n8173) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n4234), .CK(CLK), .Q(n8174) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n4235), .CK(CLK), .Q(n8175) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n4236), .CK(CLK), .Q(n8176) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n4237), .CK(CLK), .Q(n8177) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n4238), .CK(CLK), .Q(n8178) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n4239), .CK(CLK), .Q(n8179) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n4240), .CK(CLK), .Q(n8180) );
  DFF_X1 \REGISTERS_reg[8][63]  ( .D(n4241), .CK(CLK), .Q(n8181), .QN(n5492)
         );
  DFF_X1 \REGISTERS_reg[8][62]  ( .D(n4242), .CK(CLK), .Q(n8182), .QN(n5491)
         );
  DFF_X1 \REGISTERS_reg[8][61]  ( .D(n4243), .CK(CLK), .Q(n8183), .QN(n5490)
         );
  DFF_X1 \REGISTERS_reg[8][60]  ( .D(n4244), .CK(CLK), .Q(n8184), .QN(n5489)
         );
  DFF_X1 \REGISTERS_reg[8][59]  ( .D(n4245), .CK(CLK), .Q(n8185), .QN(n5488)
         );
  DFF_X1 \REGISTERS_reg[8][58]  ( .D(n4246), .CK(CLK), .Q(n8186), .QN(n5487)
         );
  DFF_X1 \REGISTERS_reg[8][57]  ( .D(n4247), .CK(CLK), .Q(n8187), .QN(n5486)
         );
  DFF_X1 \REGISTERS_reg[8][56]  ( .D(n4248), .CK(CLK), .Q(n8188), .QN(n5485)
         );
  DFF_X1 \REGISTERS_reg[8][55]  ( .D(n4249), .CK(CLK), .Q(n8189), .QN(n5484)
         );
  DFF_X1 \REGISTERS_reg[8][54]  ( .D(n4250), .CK(CLK), .Q(n8190), .QN(n5483)
         );
  DFF_X1 \REGISTERS_reg[8][53]  ( .D(n4251), .CK(CLK), .Q(n8191), .QN(n5482)
         );
  DFF_X1 \REGISTERS_reg[8][52]  ( .D(n4252), .CK(CLK), .Q(n8192), .QN(n5481)
         );
  DFF_X1 \REGISTERS_reg[8][51]  ( .D(n4253), .CK(CLK), .Q(n8193), .QN(n5480)
         );
  DFF_X1 \REGISTERS_reg[8][50]  ( .D(n4254), .CK(CLK), .Q(n8194), .QN(n5479)
         );
  DFF_X1 \REGISTERS_reg[8][49]  ( .D(n4255), .CK(CLK), .Q(n8195), .QN(n5478)
         );
  DFF_X1 \REGISTERS_reg[8][48]  ( .D(n4256), .CK(CLK), .Q(n8196), .QN(n5477)
         );
  DFF_X1 \REGISTERS_reg[8][47]  ( .D(n4257), .CK(CLK), .Q(n8197), .QN(n5476)
         );
  DFF_X1 \REGISTERS_reg[8][46]  ( .D(n4258), .CK(CLK), .Q(n8198), .QN(n5475)
         );
  DFF_X1 \REGISTERS_reg[8][45]  ( .D(n4259), .CK(CLK), .Q(n8199), .QN(n5474)
         );
  DFF_X1 \REGISTERS_reg[8][44]  ( .D(n4260), .CK(CLK), .Q(n8200), .QN(n5473)
         );
  DFF_X1 \REGISTERS_reg[8][43]  ( .D(n4261), .CK(CLK), .Q(n8201), .QN(n5472)
         );
  DFF_X1 \REGISTERS_reg[8][42]  ( .D(n4262), .CK(CLK), .Q(n8202), .QN(n5471)
         );
  DFF_X1 \REGISTERS_reg[8][41]  ( .D(n4263), .CK(CLK), .Q(n8203), .QN(n5470)
         );
  DFF_X1 \REGISTERS_reg[8][40]  ( .D(n4264), .CK(CLK), .Q(n8204), .QN(n5469)
         );
  DFF_X1 \REGISTERS_reg[8][39]  ( .D(n4265), .CK(CLK), .Q(n8205), .QN(n5468)
         );
  DFF_X1 \REGISTERS_reg[8][38]  ( .D(n4266), .CK(CLK), .Q(n8206), .QN(n5467)
         );
  DFF_X1 \REGISTERS_reg[8][37]  ( .D(n4267), .CK(CLK), .Q(n8207), .QN(n5466)
         );
  DFF_X1 \REGISTERS_reg[8][36]  ( .D(n4268), .CK(CLK), .Q(n8208), .QN(n5465)
         );
  DFF_X1 \REGISTERS_reg[8][35]  ( .D(n4269), .CK(CLK), .Q(n8209), .QN(n5464)
         );
  DFF_X1 \REGISTERS_reg[8][34]  ( .D(n4270), .CK(CLK), .Q(n8210), .QN(n5463)
         );
  DFF_X1 \REGISTERS_reg[8][33]  ( .D(n4271), .CK(CLK), .Q(n8211), .QN(n5462)
         );
  DFF_X1 \REGISTERS_reg[8][32]  ( .D(n4272), .CK(CLK), .Q(n8212), .QN(n5461)
         );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n4273), .CK(CLK), .Q(n8213), .QN(n5460)
         );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n4274), .CK(CLK), .Q(n8214), .QN(n5459)
         );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n4275), .CK(CLK), .Q(n8215), .QN(n5458)
         );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n4276), .CK(CLK), .Q(n8216), .QN(n5457)
         );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n4277), .CK(CLK), .Q(n8217), .QN(n5456)
         );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n4278), .CK(CLK), .Q(n8218), .QN(n5455)
         );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n4279), .CK(CLK), .Q(n8219), .QN(n5454)
         );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n4280), .CK(CLK), .Q(n8220), .QN(n5453)
         );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n4281), .CK(CLK), .Q(n8221), .QN(n5452)
         );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n4282), .CK(CLK), .Q(n8222), .QN(n5451)
         );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n4283), .CK(CLK), .Q(n8223), .QN(n5450)
         );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n4284), .CK(CLK), .Q(n8224), .QN(n5449)
         );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n4285), .CK(CLK), .Q(n8225), .QN(n5448)
         );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n4286), .CK(CLK), .Q(n8226), .QN(n5447)
         );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n4287), .CK(CLK), .Q(n8227), .QN(n5446)
         );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n4288), .CK(CLK), .Q(n8228), .QN(n5445)
         );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n4289), .CK(CLK), .Q(n8229), .QN(n5444)
         );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n4290), .CK(CLK), .Q(n8230), .QN(n5443)
         );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n4291), .CK(CLK), .Q(n8231), .QN(n5442)
         );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n4292), .CK(CLK), .Q(n8232), .QN(n5441)
         );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n4293), .CK(CLK), .Q(n8233), .QN(n5440)
         );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n4294), .CK(CLK), .Q(n8234), .QN(n5439)
         );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n4295), .CK(CLK), .Q(n8235), .QN(n5438) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n4296), .CK(CLK), .Q(n8236), .QN(n5437) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n4297), .CK(CLK), .Q(n8237), .QN(n5436) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n4298), .CK(CLK), .Q(n8238), .QN(n5435) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n4299), .CK(CLK), .Q(n8239), .QN(n5434) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n4300), .CK(CLK), .Q(n8240), .QN(n5433) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n4301), .CK(CLK), .Q(n8241), .QN(n5432) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n4302), .CK(CLK), .Q(n8242), .QN(n5431) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n4303), .CK(CLK), .Q(n8243), .QN(n5430) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n4304), .CK(CLK), .Q(n8244), .QN(n5429) );
  DFF_X1 \REGISTERS_reg[9][63]  ( .D(n4305), .CK(CLK), .Q(n5686), .QN(n738) );
  DFF_X1 \REGISTERS_reg[9][62]  ( .D(n4306), .CK(CLK), .Q(n5685), .QN(n739) );
  DFF_X1 \REGISTERS_reg[9][61]  ( .D(n4307), .CK(CLK), .Q(n5684), .QN(n740) );
  DFF_X1 \REGISTERS_reg[9][60]  ( .D(n4308), .CK(CLK), .Q(n5683), .QN(n741) );
  DFF_X1 \REGISTERS_reg[9][59]  ( .D(n4309), .CK(CLK), .Q(n5682), .QN(n742) );
  DFF_X1 \REGISTERS_reg[9][58]  ( .D(n4310), .CK(CLK), .Q(n5681), .QN(n743) );
  DFF_X1 \REGISTERS_reg[9][57]  ( .D(n4311), .CK(CLK), .Q(n5680), .QN(n744) );
  DFF_X1 \REGISTERS_reg[9][56]  ( .D(n4312), .CK(CLK), .Q(n5679), .QN(n745) );
  DFF_X1 \REGISTERS_reg[9][55]  ( .D(n4313), .CK(CLK), .Q(n5678), .QN(n746) );
  DFF_X1 \REGISTERS_reg[9][54]  ( .D(n4314), .CK(CLK), .Q(n5677), .QN(n747) );
  DFF_X1 \REGISTERS_reg[9][53]  ( .D(n4315), .CK(CLK), .Q(n5676), .QN(n748) );
  DFF_X1 \REGISTERS_reg[9][52]  ( .D(n4316), .CK(CLK), .Q(n5675), .QN(n749) );
  DFF_X1 \REGISTERS_reg[9][51]  ( .D(n4317), .CK(CLK), .Q(n5674), .QN(n750) );
  DFF_X1 \REGISTERS_reg[9][50]  ( .D(n4318), .CK(CLK), .Q(n5673), .QN(n751) );
  DFF_X1 \REGISTERS_reg[9][49]  ( .D(n4319), .CK(CLK), .Q(n5672), .QN(n752) );
  DFF_X1 \REGISTERS_reg[9][48]  ( .D(n4320), .CK(CLK), .Q(n5671), .QN(n753) );
  DFF_X1 \REGISTERS_reg[9][47]  ( .D(n4321), .CK(CLK), .Q(n5670), .QN(n754) );
  DFF_X1 \REGISTERS_reg[9][46]  ( .D(n4322), .CK(CLK), .Q(n5669), .QN(n755) );
  DFF_X1 \REGISTERS_reg[9][45]  ( .D(n4323), .CK(CLK), .Q(n5668), .QN(n756) );
  DFF_X1 \REGISTERS_reg[9][44]  ( .D(n4324), .CK(CLK), .Q(n5667), .QN(n757) );
  DFF_X1 \REGISTERS_reg[9][43]  ( .D(n4325), .CK(CLK), .Q(n5666), .QN(n758) );
  DFF_X1 \REGISTERS_reg[9][42]  ( .D(n4326), .CK(CLK), .Q(n5665), .QN(n759) );
  DFF_X1 \REGISTERS_reg[9][41]  ( .D(n4327), .CK(CLK), .Q(n5664), .QN(n760) );
  DFF_X1 \REGISTERS_reg[9][40]  ( .D(n4328), .CK(CLK), .Q(n5663), .QN(n761) );
  DFF_X1 \REGISTERS_reg[9][39]  ( .D(n4329), .CK(CLK), .Q(n5662), .QN(n762) );
  DFF_X1 \REGISTERS_reg[9][38]  ( .D(n4330), .CK(CLK), .Q(n5661), .QN(n763) );
  DFF_X1 \REGISTERS_reg[9][37]  ( .D(n4331), .CK(CLK), .Q(n5660), .QN(n764) );
  DFF_X1 \REGISTERS_reg[9][36]  ( .D(n4332), .CK(CLK), .Q(n5659), .QN(n765) );
  DFF_X1 \REGISTERS_reg[9][35]  ( .D(n4333), .CK(CLK), .Q(n5658), .QN(n766) );
  DFF_X1 \REGISTERS_reg[9][34]  ( .D(n4334), .CK(CLK), .Q(n5657), .QN(n767) );
  DFF_X1 \REGISTERS_reg[9][33]  ( .D(n4335), .CK(CLK), .Q(n5656), .QN(n768) );
  DFF_X1 \REGISTERS_reg[9][32]  ( .D(n4336), .CK(CLK), .Q(n5655), .QN(n769) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n4337), .CK(CLK), .Q(n5654), .QN(n770) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n4338), .CK(CLK), .Q(n5653), .QN(n771) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n4339), .CK(CLK), .Q(n5652), .QN(n772) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n4340), .CK(CLK), .Q(n5651), .QN(n773) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n4341), .CK(CLK), .Q(n5650), .QN(n774) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n4342), .CK(CLK), .Q(n5649), .QN(n775) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n4343), .CK(CLK), .Q(n5648), .QN(n776) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n4344), .CK(CLK), .Q(n5647), .QN(n777) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n4345), .CK(CLK), .Q(n5646), .QN(n778) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n4346), .CK(CLK), .Q(n5645), .QN(n779) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n4347), .CK(CLK), .Q(n5644), .QN(n780) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n4348), .CK(CLK), .Q(n5643), .QN(n781) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n4349), .CK(CLK), .Q(n5642), .QN(n782) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n4350), .CK(CLK), .Q(n5641), .QN(n783) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n4351), .CK(CLK), .Q(n5640), .QN(n784) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n4352), .CK(CLK), .Q(n5639), .QN(n785) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n4353), .CK(CLK), .Q(n5638), .QN(n786) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n4354), .CK(CLK), .Q(n5637), .QN(n787) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n4355), .CK(CLK), .Q(n5636), .QN(n788) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n4356), .CK(CLK), .Q(n5635), .QN(n789) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n4357), .CK(CLK), .Q(n5634), .QN(n790) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n4358), .CK(CLK), .Q(n5633), .QN(n791) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n4359), .CK(CLK), .Q(n5632), .QN(n792) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n4360), .CK(CLK), .Q(n5631), .QN(n793) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n4361), .CK(CLK), .Q(n5630), .QN(n794) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n4362), .CK(CLK), .Q(n5629), .QN(n795) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n4363), .CK(CLK), .Q(n5628), .QN(n796) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n4364), .CK(CLK), .Q(n5627), .QN(n797) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n4365), .CK(CLK), .Q(n5626), .QN(n798) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n4366), .CK(CLK), .Q(n5625), .QN(n799) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n4367), .CK(CLK), .Q(n5624), .QN(n800) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n4368), .CK(CLK), .Q(n5623), .QN(n801) );
  DFF_X1 \REGISTERS_reg[10][63]  ( .D(n4369), .CK(CLK), .Q(n5364), .QN(n802)
         );
  DFF_X1 \REGISTERS_reg[10][62]  ( .D(n4370), .CK(CLK), .Q(n5363), .QN(n803)
         );
  DFF_X1 \REGISTERS_reg[10][61]  ( .D(n4371), .CK(CLK), .Q(n5362), .QN(n804)
         );
  DFF_X1 \REGISTERS_reg[10][60]  ( .D(n4372), .CK(CLK), .Q(n5361), .QN(n805)
         );
  DFF_X1 \REGISTERS_reg[10][59]  ( .D(n4373), .CK(CLK), .Q(n5360), .QN(n806)
         );
  DFF_X1 \REGISTERS_reg[10][58]  ( .D(n4374), .CK(CLK), .Q(n5359), .QN(n807)
         );
  DFF_X1 \REGISTERS_reg[10][57]  ( .D(n4375), .CK(CLK), .Q(n5358), .QN(n808)
         );
  DFF_X1 \REGISTERS_reg[10][56]  ( .D(n4376), .CK(CLK), .Q(n5357), .QN(n809)
         );
  DFF_X1 \REGISTERS_reg[10][55]  ( .D(n4377), .CK(CLK), .Q(n5356), .QN(n810)
         );
  DFF_X1 \REGISTERS_reg[10][54]  ( .D(n4378), .CK(CLK), .Q(n5355), .QN(n811)
         );
  DFF_X1 \REGISTERS_reg[10][53]  ( .D(n4379), .CK(CLK), .Q(n5354), .QN(n812)
         );
  DFF_X1 \REGISTERS_reg[10][52]  ( .D(n4380), .CK(CLK), .Q(n5353), .QN(n813)
         );
  DFF_X1 \REGISTERS_reg[10][51]  ( .D(n4381), .CK(CLK), .Q(n5352), .QN(n814)
         );
  DFF_X1 \REGISTERS_reg[10][50]  ( .D(n4382), .CK(CLK), .Q(n5351), .QN(n815)
         );
  DFF_X1 \REGISTERS_reg[10][49]  ( .D(n4383), .CK(CLK), .Q(n5350), .QN(n816)
         );
  DFF_X1 \REGISTERS_reg[10][48]  ( .D(n4384), .CK(CLK), .Q(n5349), .QN(n817)
         );
  DFF_X1 \REGISTERS_reg[10][47]  ( .D(n4385), .CK(CLK), .Q(n5348), .QN(n818)
         );
  DFF_X1 \REGISTERS_reg[10][46]  ( .D(n4386), .CK(CLK), .Q(n5347), .QN(n819)
         );
  DFF_X1 \REGISTERS_reg[10][45]  ( .D(n4387), .CK(CLK), .Q(n5346), .QN(n820)
         );
  DFF_X1 \REGISTERS_reg[10][44]  ( .D(n4388), .CK(CLK), .Q(n5345), .QN(n821)
         );
  DFF_X1 \REGISTERS_reg[10][43]  ( .D(n4389), .CK(CLK), .Q(n5344), .QN(n822)
         );
  DFF_X1 \REGISTERS_reg[10][42]  ( .D(n4390), .CK(CLK), .Q(n5343), .QN(n823)
         );
  DFF_X1 \REGISTERS_reg[10][41]  ( .D(n4391), .CK(CLK), .Q(n5342), .QN(n824)
         );
  DFF_X1 \REGISTERS_reg[10][40]  ( .D(n4392), .CK(CLK), .Q(n5341), .QN(n825)
         );
  DFF_X1 \REGISTERS_reg[10][39]  ( .D(n4393), .CK(CLK), .Q(n5340), .QN(n826)
         );
  DFF_X1 \REGISTERS_reg[10][38]  ( .D(n4394), .CK(CLK), .Q(n5339), .QN(n827)
         );
  DFF_X1 \REGISTERS_reg[10][37]  ( .D(n4395), .CK(CLK), .Q(n5338), .QN(n828)
         );
  DFF_X1 \REGISTERS_reg[10][36]  ( .D(n4396), .CK(CLK), .Q(n5337), .QN(n829)
         );
  DFF_X1 \REGISTERS_reg[10][35]  ( .D(n4397), .CK(CLK), .Q(n5336), .QN(n830)
         );
  DFF_X1 \REGISTERS_reg[10][34]  ( .D(n4398), .CK(CLK), .Q(n5335), .QN(n831)
         );
  DFF_X1 \REGISTERS_reg[10][33]  ( .D(n4399), .CK(CLK), .Q(n5334), .QN(n832)
         );
  DFF_X1 \REGISTERS_reg[10][32]  ( .D(n4400), .CK(CLK), .Q(n5333), .QN(n833)
         );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n4401), .CK(CLK), .Q(n5332), .QN(n834)
         );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n4402), .CK(CLK), .Q(n5331), .QN(n835)
         );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n4403), .CK(CLK), .Q(n5330), .QN(n836)
         );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n4404), .CK(CLK), .Q(n5329), .QN(n837)
         );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n4405), .CK(CLK), .Q(n5328), .QN(n838)
         );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n4406), .CK(CLK), .Q(n5327), .QN(n839)
         );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n4407), .CK(CLK), .Q(n5326), .QN(n840)
         );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n4408), .CK(CLK), .Q(n5325), .QN(n841)
         );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n4409), .CK(CLK), .Q(n5324), .QN(n842)
         );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n4410), .CK(CLK), .Q(n5323), .QN(n843)
         );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n4411), .CK(CLK), .Q(n5322), .QN(n844)
         );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n4412), .CK(CLK), .Q(n5321), .QN(n845)
         );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n4413), .CK(CLK), .Q(n5320), .QN(n846)
         );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n4414), .CK(CLK), .Q(n5319), .QN(n847)
         );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n4415), .CK(CLK), .Q(n5318), .QN(n848)
         );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n4416), .CK(CLK), .Q(n5317), .QN(n849)
         );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n4417), .CK(CLK), .Q(n5316), .QN(n850)
         );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n4418), .CK(CLK), .Q(n5315), .QN(n851)
         );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n4419), .CK(CLK), .Q(n5314), .QN(n852)
         );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n4420), .CK(CLK), .Q(n5313), .QN(n853)
         );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n4421), .CK(CLK), .Q(n5312), .QN(n854)
         );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n4422), .CK(CLK), .Q(n5311), .QN(n855)
         );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n4423), .CK(CLK), .Q(n5310), .QN(n856) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n4424), .CK(CLK), .Q(n5309), .QN(n857) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n4425), .CK(CLK), .Q(n5308), .QN(n858) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n4426), .CK(CLK), .Q(n5307), .QN(n859) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n4427), .CK(CLK), .Q(n5306), .QN(n860) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n4428), .CK(CLK), .Q(n5305), .QN(n861) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n4429), .CK(CLK), .Q(n5304), .QN(n862) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n4430), .CK(CLK), .Q(n5303), .QN(n863) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n4431), .CK(CLK), .Q(n5302), .QN(n864) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n4432), .CK(CLK), .Q(n5301), .QN(n865) );
  DFF_X1 \REGISTERS_reg[11][63]  ( .D(n4433), .CK(CLK), .Q(n5153), .QN(n866)
         );
  DFF_X1 \REGISTERS_reg[11][62]  ( .D(n4434), .CK(CLK), .Q(n5152), .QN(n867)
         );
  DFF_X1 \REGISTERS_reg[11][61]  ( .D(n4435), .CK(CLK), .Q(n5151), .QN(n868)
         );
  DFF_X1 \REGISTERS_reg[11][60]  ( .D(n4436), .CK(CLK), .Q(n5150), .QN(n869)
         );
  DFF_X1 \REGISTERS_reg[11][59]  ( .D(n4437), .CK(CLK), .Q(n5149), .QN(n870)
         );
  DFF_X1 \REGISTERS_reg[11][58]  ( .D(n4438), .CK(CLK), .Q(n5148), .QN(n871)
         );
  DFF_X1 \REGISTERS_reg[11][57]  ( .D(n4439), .CK(CLK), .Q(n5147), .QN(n872)
         );
  DFF_X1 \REGISTERS_reg[11][56]  ( .D(n4440), .CK(CLK), .Q(n5146), .QN(n873)
         );
  DFF_X1 \REGISTERS_reg[11][55]  ( .D(n4441), .CK(CLK), .Q(n5145), .QN(n874)
         );
  DFF_X1 \REGISTERS_reg[11][54]  ( .D(n4442), .CK(CLK), .Q(n5144), .QN(n875)
         );
  DFF_X1 \REGISTERS_reg[11][53]  ( .D(n4443), .CK(CLK), .Q(n5143), .QN(n876)
         );
  DFF_X1 \REGISTERS_reg[11][52]  ( .D(n4444), .CK(CLK), .Q(n5142), .QN(n877)
         );
  DFF_X1 \REGISTERS_reg[11][51]  ( .D(n4445), .CK(CLK), .Q(n5141), .QN(n878)
         );
  DFF_X1 \REGISTERS_reg[11][50]  ( .D(n4446), .CK(CLK), .Q(n5140), .QN(n879)
         );
  DFF_X1 \REGISTERS_reg[11][49]  ( .D(n4447), .CK(CLK), .Q(n5139), .QN(n880)
         );
  DFF_X1 \REGISTERS_reg[11][48]  ( .D(n4448), .CK(CLK), .Q(n5138), .QN(n881)
         );
  DFF_X1 \REGISTERS_reg[11][47]  ( .D(n4449), .CK(CLK), .Q(n5137), .QN(n882)
         );
  DFF_X1 \REGISTERS_reg[11][46]  ( .D(n4450), .CK(CLK), .Q(n5136), .QN(n883)
         );
  DFF_X1 \REGISTERS_reg[11][45]  ( .D(n4451), .CK(CLK), .Q(n5135), .QN(n884)
         );
  DFF_X1 \REGISTERS_reg[11][44]  ( .D(n4452), .CK(CLK), .Q(n5134), .QN(n885)
         );
  DFF_X1 \REGISTERS_reg[11][43]  ( .D(n4453), .CK(CLK), .Q(n5133), .QN(n886)
         );
  DFF_X1 \REGISTERS_reg[11][42]  ( .D(n4454), .CK(CLK), .Q(n5132), .QN(n887)
         );
  DFF_X1 \REGISTERS_reg[11][41]  ( .D(n4455), .CK(CLK), .Q(n5131), .QN(n888)
         );
  DFF_X1 \REGISTERS_reg[11][40]  ( .D(n4456), .CK(CLK), .Q(n5130), .QN(n889)
         );
  DFF_X1 \REGISTERS_reg[11][39]  ( .D(n4457), .CK(CLK), .Q(n5129), .QN(n890)
         );
  DFF_X1 \REGISTERS_reg[11][38]  ( .D(n4458), .CK(CLK), .Q(n5128), .QN(n891)
         );
  DFF_X1 \REGISTERS_reg[11][37]  ( .D(n4459), .CK(CLK), .Q(n5127), .QN(n892)
         );
  DFF_X1 \REGISTERS_reg[11][36]  ( .D(n4460), .CK(CLK), .Q(n5126), .QN(n893)
         );
  DFF_X1 \REGISTERS_reg[11][35]  ( .D(n4461), .CK(CLK), .Q(n5125), .QN(n894)
         );
  DFF_X1 \REGISTERS_reg[11][34]  ( .D(n4462), .CK(CLK), .Q(n5124), .QN(n895)
         );
  DFF_X1 \REGISTERS_reg[11][33]  ( .D(n4463), .CK(CLK), .Q(n5123), .QN(n896)
         );
  DFF_X1 \REGISTERS_reg[11][32]  ( .D(n4464), .CK(CLK), .Q(n5122), .QN(n897)
         );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n4465), .CK(CLK), .Q(n5121), .QN(n898)
         );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n4466), .CK(CLK), .Q(n5120), .QN(n899)
         );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n4467), .CK(CLK), .Q(n5119), .QN(n900)
         );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n4468), .CK(CLK), .Q(n5118), .QN(n901)
         );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n4469), .CK(CLK), .Q(n5117), .QN(n902)
         );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n4470), .CK(CLK), .Q(n5116), .QN(n903)
         );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n4471), .CK(CLK), .Q(n5115), .QN(n904)
         );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n4472), .CK(CLK), .Q(n5114), .QN(n905)
         );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n4473), .CK(CLK), .Q(n5113), .QN(n906)
         );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n4474), .CK(CLK), .Q(n5112), .QN(n907)
         );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n4475), .CK(CLK), .Q(n5111), .QN(n908)
         );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n4476), .CK(CLK), .Q(n5110), .QN(n909)
         );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n4477), .CK(CLK), .Q(n5109), .QN(n910)
         );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n4478), .CK(CLK), .Q(n5108), .QN(n911)
         );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n4479), .CK(CLK), .Q(n5107), .QN(n912)
         );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n4480), .CK(CLK), .Q(n5106), .QN(n913)
         );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n4481), .CK(CLK), .Q(n5105), .QN(n914)
         );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n4482), .CK(CLK), .Q(n5104), .QN(n915)
         );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n4483), .CK(CLK), .Q(n5103), .QN(n916)
         );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n4484), .CK(CLK), .Q(n5102), .QN(n917)
         );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n4485), .CK(CLK), .Q(n5101), .QN(n918)
         );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n4486), .CK(CLK), .Q(n5100), .QN(n919)
         );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n4487), .CK(CLK), .Q(n5099), .QN(n920) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n4488), .CK(CLK), .Q(n5098), .QN(n921) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n4489), .CK(CLK), .Q(n5097), .QN(n922) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n4490), .CK(CLK), .Q(n5096), .QN(n923) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n4491), .CK(CLK), .Q(n5095), .QN(n924) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n4492), .CK(CLK), .Q(n5094), .QN(n925) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n4493), .CK(CLK), .Q(n5093), .QN(n926) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n4494), .CK(CLK), .Q(n5092), .QN(n927) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n4495), .CK(CLK), .Q(n5091), .QN(n928) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n4496), .CK(CLK), .Q(n5090), .QN(n929) );
  DFF_X1 \REGISTERS_reg[12][63]  ( .D(n4497), .CK(CLK), .Q(n5750), .QN(n930)
         );
  DFF_X1 \REGISTERS_reg[12][62]  ( .D(n4498), .CK(CLK), .Q(n5749), .QN(n931)
         );
  DFF_X1 \REGISTERS_reg[12][61]  ( .D(n4499), .CK(CLK), .Q(n5748), .QN(n932)
         );
  DFF_X1 \REGISTERS_reg[12][60]  ( .D(n4500), .CK(CLK), .Q(n5747), .QN(n933)
         );
  DFF_X1 \REGISTERS_reg[12][59]  ( .D(n4501), .CK(CLK), .Q(n5746), .QN(n934)
         );
  DFF_X1 \REGISTERS_reg[12][58]  ( .D(n4502), .CK(CLK), .Q(n5745), .QN(n935)
         );
  DFF_X1 \REGISTERS_reg[12][57]  ( .D(n4503), .CK(CLK), .Q(n5744), .QN(n936)
         );
  DFF_X1 \REGISTERS_reg[12][56]  ( .D(n4504), .CK(CLK), .Q(n5743), .QN(n937)
         );
  DFF_X1 \REGISTERS_reg[12][55]  ( .D(n4505), .CK(CLK), .Q(n5742), .QN(n938)
         );
  DFF_X1 \REGISTERS_reg[12][54]  ( .D(n4506), .CK(CLK), .Q(n5741), .QN(n939)
         );
  DFF_X1 \REGISTERS_reg[12][53]  ( .D(n4507), .CK(CLK), .Q(n5740), .QN(n940)
         );
  DFF_X1 \REGISTERS_reg[12][52]  ( .D(n4508), .CK(CLK), .Q(n5739), .QN(n941)
         );
  DFF_X1 \REGISTERS_reg[12][51]  ( .D(n4509), .CK(CLK), .Q(n5738), .QN(n942)
         );
  DFF_X1 \REGISTERS_reg[12][50]  ( .D(n4510), .CK(CLK), .Q(n5737), .QN(n943)
         );
  DFF_X1 \REGISTERS_reg[12][49]  ( .D(n4511), .CK(CLK), .Q(n5736), .QN(n944)
         );
  DFF_X1 \REGISTERS_reg[12][48]  ( .D(n4512), .CK(CLK), .Q(n5735), .QN(n945)
         );
  DFF_X1 \REGISTERS_reg[12][47]  ( .D(n4513), .CK(CLK), .Q(n5734), .QN(n946)
         );
  DFF_X1 \REGISTERS_reg[12][46]  ( .D(n4514), .CK(CLK), .Q(n5733), .QN(n947)
         );
  DFF_X1 \REGISTERS_reg[12][45]  ( .D(n4515), .CK(CLK), .Q(n5732), .QN(n948)
         );
  DFF_X1 \REGISTERS_reg[12][44]  ( .D(n4516), .CK(CLK), .Q(n5731), .QN(n949)
         );
  DFF_X1 \REGISTERS_reg[12][43]  ( .D(n4517), .CK(CLK), .Q(n5730), .QN(n950)
         );
  DFF_X1 \REGISTERS_reg[12][42]  ( .D(n4518), .CK(CLK), .Q(n5729), .QN(n951)
         );
  DFF_X1 \REGISTERS_reg[12][41]  ( .D(n4519), .CK(CLK), .Q(n5728), .QN(n952)
         );
  DFF_X1 \REGISTERS_reg[12][40]  ( .D(n4520), .CK(CLK), .Q(n5727), .QN(n953)
         );
  DFF_X1 \REGISTERS_reg[12][39]  ( .D(n4521), .CK(CLK), .Q(n5726), .QN(n954)
         );
  DFF_X1 \REGISTERS_reg[12][38]  ( .D(n4522), .CK(CLK), .Q(n5725), .QN(n955)
         );
  DFF_X1 \REGISTERS_reg[12][37]  ( .D(n4523), .CK(CLK), .Q(n5724), .QN(n956)
         );
  DFF_X1 \REGISTERS_reg[12][36]  ( .D(n4524), .CK(CLK), .Q(n5723), .QN(n957)
         );
  DFF_X1 \REGISTERS_reg[12][35]  ( .D(n4525), .CK(CLK), .Q(n5722), .QN(n958)
         );
  DFF_X1 \REGISTERS_reg[12][34]  ( .D(n4526), .CK(CLK), .Q(n5721), .QN(n959)
         );
  DFF_X1 \REGISTERS_reg[12][33]  ( .D(n4527), .CK(CLK), .Q(n5720), .QN(n960)
         );
  DFF_X1 \REGISTERS_reg[12][32]  ( .D(n4528), .CK(CLK), .Q(n5719), .QN(n961)
         );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n4529), .CK(CLK), .Q(n5718), .QN(n962)
         );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n4530), .CK(CLK), .Q(n5717), .QN(n963)
         );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n4531), .CK(CLK), .Q(n5716), .QN(n964)
         );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n4532), .CK(CLK), .Q(n5715), .QN(n965)
         );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n4533), .CK(CLK), .Q(n5714), .QN(n966)
         );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n4534), .CK(CLK), .Q(n5713), .QN(n967)
         );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n4535), .CK(CLK), .Q(n5712), .QN(n968)
         );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n4536), .CK(CLK), .Q(n5711), .QN(n969)
         );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n4537), .CK(CLK), .Q(n5710), .QN(n970)
         );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n4538), .CK(CLK), .Q(n5709), .QN(n971)
         );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n4539), .CK(CLK), .Q(n5708), .QN(n972)
         );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n4540), .CK(CLK), .Q(n5707), .QN(n973)
         );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n4541), .CK(CLK), .Q(n5706), .QN(n974)
         );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n4542), .CK(CLK), .Q(n5705), .QN(n975)
         );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n4543), .CK(CLK), .Q(n5704), .QN(n976)
         );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n4544), .CK(CLK), .Q(n5703), .QN(n977)
         );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n4545), .CK(CLK), .Q(n5702), .QN(n978)
         );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n4546), .CK(CLK), .Q(n5701), .QN(n979)
         );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n4547), .CK(CLK), .Q(n5700), .QN(n980)
         );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n4548), .CK(CLK), .Q(n5699), .QN(n981)
         );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n4549), .CK(CLK), .Q(n5698), .QN(n982)
         );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n4550), .CK(CLK), .Q(n5697), .QN(n983)
         );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n4551), .CK(CLK), .Q(n5696), .QN(n984) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n4552), .CK(CLK), .Q(n5695), .QN(n985) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n4553), .CK(CLK), .Q(n5694), .QN(n986) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n4554), .CK(CLK), .Q(n5693), .QN(n987) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n4555), .CK(CLK), .Q(n5692), .QN(n988) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n4556), .CK(CLK), .Q(n5691), .QN(n989) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n4557), .CK(CLK), .Q(n5690), .QN(n990) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n4558), .CK(CLK), .Q(n5689), .QN(n991) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n4559), .CK(CLK), .Q(n5688), .QN(n992) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n4560), .CK(CLK), .Q(n5687), .QN(n993) );
  DFF_X1 \REGISTERS_reg[13][63]  ( .D(n4561), .CK(CLK), .Q(n5217), .QN(n994)
         );
  DFF_X1 \REGISTERS_reg[13][62]  ( .D(n4562), .CK(CLK), .Q(n5216), .QN(n995)
         );
  DFF_X1 \REGISTERS_reg[13][61]  ( .D(n4563), .CK(CLK), .Q(n5215), .QN(n996)
         );
  DFF_X1 \REGISTERS_reg[13][60]  ( .D(n4564), .CK(CLK), .Q(n5214), .QN(n997)
         );
  DFF_X1 \REGISTERS_reg[13][59]  ( .D(n4565), .CK(CLK), .Q(n5213), .QN(n998)
         );
  DFF_X1 \REGISTERS_reg[13][58]  ( .D(n4566), .CK(CLK), .Q(n5212), .QN(n999)
         );
  DFF_X1 \REGISTERS_reg[13][57]  ( .D(n4567), .CK(CLK), .Q(n5211), .QN(n1000)
         );
  DFF_X1 \REGISTERS_reg[13][56]  ( .D(n4568), .CK(CLK), .Q(n5210), .QN(n1001)
         );
  DFF_X1 \REGISTERS_reg[13][55]  ( .D(n4569), .CK(CLK), .Q(n5209), .QN(n1002)
         );
  DFF_X1 \REGISTERS_reg[13][54]  ( .D(n4570), .CK(CLK), .Q(n5208), .QN(n1003)
         );
  DFF_X1 \REGISTERS_reg[13][53]  ( .D(n4571), .CK(CLK), .Q(n5207), .QN(n1004)
         );
  DFF_X1 \REGISTERS_reg[13][52]  ( .D(n4572), .CK(CLK), .Q(n5206), .QN(n1005)
         );
  DFF_X1 \REGISTERS_reg[13][51]  ( .D(n4573), .CK(CLK), .Q(n5205), .QN(n1006)
         );
  DFF_X1 \REGISTERS_reg[13][50]  ( .D(n4574), .CK(CLK), .Q(n5204), .QN(n1007)
         );
  DFF_X1 \REGISTERS_reg[13][49]  ( .D(n4575), .CK(CLK), .Q(n5203), .QN(n1008)
         );
  DFF_X1 \REGISTERS_reg[13][48]  ( .D(n4576), .CK(CLK), .Q(n5202), .QN(n1009)
         );
  DFF_X1 \REGISTERS_reg[13][47]  ( .D(n4577), .CK(CLK), .Q(n5201), .QN(n1010)
         );
  DFF_X1 \REGISTERS_reg[13][46]  ( .D(n4578), .CK(CLK), .Q(n5200), .QN(n1011)
         );
  DFF_X1 \REGISTERS_reg[13][45]  ( .D(n4579), .CK(CLK), .Q(n5199), .QN(n1012)
         );
  DFF_X1 \REGISTERS_reg[13][44]  ( .D(n4580), .CK(CLK), .Q(n5198), .QN(n1013)
         );
  DFF_X1 \REGISTERS_reg[13][43]  ( .D(n4581), .CK(CLK), .Q(n5197), .QN(n1014)
         );
  DFF_X1 \REGISTERS_reg[13][42]  ( .D(n4582), .CK(CLK), .Q(n5196), .QN(n1015)
         );
  DFF_X1 \REGISTERS_reg[13][41]  ( .D(n4583), .CK(CLK), .Q(n5195), .QN(n1016)
         );
  DFF_X1 \REGISTERS_reg[13][40]  ( .D(n4584), .CK(CLK), .Q(n5194), .QN(n1017)
         );
  DFF_X1 \REGISTERS_reg[13][39]  ( .D(n4585), .CK(CLK), .Q(n5193), .QN(n1018)
         );
  DFF_X1 \REGISTERS_reg[13][38]  ( .D(n4586), .CK(CLK), .Q(n5192), .QN(n1019)
         );
  DFF_X1 \REGISTERS_reg[13][37]  ( .D(n4587), .CK(CLK), .Q(n5191), .QN(n1020)
         );
  DFF_X1 \REGISTERS_reg[13][36]  ( .D(n4588), .CK(CLK), .Q(n5190), .QN(n1021)
         );
  DFF_X1 \REGISTERS_reg[13][35]  ( .D(n4589), .CK(CLK), .Q(n5189), .QN(n1022)
         );
  DFF_X1 \REGISTERS_reg[13][34]  ( .D(n4590), .CK(CLK), .Q(n5188), .QN(n1023)
         );
  DFF_X1 \REGISTERS_reg[13][33]  ( .D(n4591), .CK(CLK), .Q(n5187), .QN(n1024)
         );
  DFF_X1 \REGISTERS_reg[13][32]  ( .D(n4592), .CK(CLK), .Q(n5186), .QN(n1025)
         );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n4593), .CK(CLK), .Q(n5185), .QN(n1026)
         );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n4594), .CK(CLK), .Q(n5184), .QN(n1027)
         );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n4595), .CK(CLK), .Q(n5183), .QN(n1028)
         );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n4596), .CK(CLK), .Q(n5182), .QN(n1029)
         );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n4597), .CK(CLK), .Q(n5181), .QN(n1030)
         );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n4598), .CK(CLK), .Q(n5180), .QN(n1031)
         );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n4599), .CK(CLK), .Q(n5179), .QN(n1032)
         );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n4600), .CK(CLK), .Q(n5178), .QN(n1033)
         );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n4601), .CK(CLK), .Q(n5177), .QN(n1034)
         );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n4602), .CK(CLK), .Q(n5176), .QN(n1035)
         );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n4603), .CK(CLK), .Q(n5175), .QN(n1036)
         );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n4604), .CK(CLK), .Q(n5174), .QN(n1037)
         );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n4605), .CK(CLK), .Q(n5173), .QN(n1038)
         );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n4606), .CK(CLK), .Q(n5172), .QN(n1039)
         );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n4607), .CK(CLK), .Q(n5171), .QN(n1040)
         );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n4608), .CK(CLK), .Q(n5170), .QN(n1041)
         );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n4609), .CK(CLK), .Q(n5169), .QN(n1042)
         );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n4610), .CK(CLK), .Q(n5168), .QN(n1043)
         );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n4611), .CK(CLK), .Q(n5167), .QN(n1044)
         );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n4612), .CK(CLK), .Q(n5166), .QN(n1045)
         );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n4613), .CK(CLK), .Q(n5165), .QN(n1046)
         );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n4614), .CK(CLK), .Q(n5164), .QN(n1047)
         );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n4615), .CK(CLK), .Q(n5163), .QN(n1048)
         );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n4616), .CK(CLK), .Q(n5162), .QN(n1049)
         );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n4617), .CK(CLK), .Q(n5161), .QN(n1050)
         );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n4618), .CK(CLK), .Q(n5160), .QN(n1051)
         );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n4619), .CK(CLK), .Q(n5159), .QN(n1052)
         );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n4620), .CK(CLK), .Q(n5158), .QN(n1053)
         );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n4621), .CK(CLK), .Q(n5157), .QN(n1054)
         );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n4622), .CK(CLK), .Q(n5156), .QN(n1055)
         );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n4623), .CK(CLK), .Q(n5155), .QN(n1056)
         );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n4624), .CK(CLK), .Q(n5154), .QN(n1057)
         );
  DFF_X1 \REGISTERS_reg[14][63]  ( .D(n4625), .CK(CLK), .Q(n4958), .QN(n1058)
         );
  DFF_X1 \REGISTERS_reg[14][62]  ( .D(n4626), .CK(CLK), .Q(n4957), .QN(n1059)
         );
  DFF_X1 \REGISTERS_reg[14][61]  ( .D(n4627), .CK(CLK), .Q(n4956), .QN(n1060)
         );
  DFF_X1 \REGISTERS_reg[14][60]  ( .D(n4628), .CK(CLK), .Q(n4955), .QN(n1061)
         );
  DFF_X1 \REGISTERS_reg[14][59]  ( .D(n4629), .CK(CLK), .Q(n4954), .QN(n1062)
         );
  DFF_X1 \REGISTERS_reg[14][58]  ( .D(n4630), .CK(CLK), .Q(n4953), .QN(n1063)
         );
  DFF_X1 \REGISTERS_reg[14][57]  ( .D(n4631), .CK(CLK), .Q(n4952), .QN(n1064)
         );
  DFF_X1 \REGISTERS_reg[14][56]  ( .D(n4632), .CK(CLK), .Q(n4951), .QN(n1065)
         );
  DFF_X1 \REGISTERS_reg[14][55]  ( .D(n4633), .CK(CLK), .Q(n4950), .QN(n1066)
         );
  DFF_X1 \REGISTERS_reg[14][54]  ( .D(n4634), .CK(CLK), .Q(n4949), .QN(n1067)
         );
  DFF_X1 \REGISTERS_reg[14][53]  ( .D(n4635), .CK(CLK), .Q(n4948), .QN(n1068)
         );
  DFF_X1 \REGISTERS_reg[14][52]  ( .D(n4636), .CK(CLK), .Q(n4947), .QN(n1069)
         );
  DFF_X1 \REGISTERS_reg[14][51]  ( .D(n4637), .CK(CLK), .Q(n4946), .QN(n1070)
         );
  DFF_X1 \REGISTERS_reg[14][50]  ( .D(n4638), .CK(CLK), .Q(n4945), .QN(n1071)
         );
  DFF_X1 \REGISTERS_reg[14][49]  ( .D(n4639), .CK(CLK), .Q(n4944), .QN(n1072)
         );
  DFF_X1 \REGISTERS_reg[14][48]  ( .D(n4640), .CK(CLK), .Q(n4943), .QN(n1073)
         );
  DFF_X1 \REGISTERS_reg[14][47]  ( .D(n4641), .CK(CLK), .Q(n4942), .QN(n1074)
         );
  DFF_X1 \REGISTERS_reg[14][46]  ( .D(n4642), .CK(CLK), .Q(n4941), .QN(n1075)
         );
  DFF_X1 \REGISTERS_reg[14][45]  ( .D(n4643), .CK(CLK), .Q(n4940), .QN(n1076)
         );
  DFF_X1 \REGISTERS_reg[14][44]  ( .D(n4644), .CK(CLK), .Q(n4939), .QN(n1077)
         );
  DFF_X1 \REGISTERS_reg[14][43]  ( .D(n4645), .CK(CLK), .Q(n4938), .QN(n1078)
         );
  DFF_X1 \REGISTERS_reg[14][42]  ( .D(n4646), .CK(CLK), .Q(n4937), .QN(n1079)
         );
  DFF_X1 \REGISTERS_reg[14][41]  ( .D(n4647), .CK(CLK), .Q(n4936), .QN(n1080)
         );
  DFF_X1 \REGISTERS_reg[14][40]  ( .D(n4648), .CK(CLK), .Q(n4935), .QN(n1081)
         );
  DFF_X1 \REGISTERS_reg[14][39]  ( .D(n4649), .CK(CLK), .Q(n4934), .QN(n1082)
         );
  DFF_X1 \REGISTERS_reg[14][38]  ( .D(n4650), .CK(CLK), .Q(n4933), .QN(n1083)
         );
  DFF_X1 \REGISTERS_reg[14][37]  ( .D(n4651), .CK(CLK), .Q(n4932), .QN(n1084)
         );
  DFF_X1 \REGISTERS_reg[14][36]  ( .D(n4652), .CK(CLK), .Q(n4931), .QN(n1085)
         );
  DFF_X1 \REGISTERS_reg[14][35]  ( .D(n4653), .CK(CLK), .Q(n4930), .QN(n1086)
         );
  DFF_X1 \REGISTERS_reg[14][34]  ( .D(n4654), .CK(CLK), .Q(n4929), .QN(n1087)
         );
  DFF_X1 \REGISTERS_reg[14][33]  ( .D(n4655), .CK(CLK), .Q(n4928), .QN(n1088)
         );
  DFF_X1 \REGISTERS_reg[14][32]  ( .D(n4656), .CK(CLK), .Q(n4927), .QN(n1089)
         );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n4657), .CK(CLK), .Q(n4926), .QN(n1090)
         );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n4658), .CK(CLK), .Q(n4925), .QN(n1091)
         );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n4659), .CK(CLK), .Q(n4924), .QN(n1092)
         );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n4660), .CK(CLK), .Q(n4923), .QN(n1093)
         );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n4661), .CK(CLK), .Q(n4922), .QN(n1094)
         );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n4662), .CK(CLK), .Q(n4921), .QN(n1095)
         );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n4663), .CK(CLK), .Q(n4920), .QN(n1096)
         );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n4664), .CK(CLK), .Q(n4919), .QN(n1097)
         );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n4665), .CK(CLK), .Q(n4918), .QN(n1098)
         );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n4666), .CK(CLK), .Q(n4917), .QN(n1099)
         );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n4667), .CK(CLK), .Q(n4916), .QN(n1100)
         );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n4668), .CK(CLK), .Q(n4915), .QN(n1101)
         );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n4669), .CK(CLK), .Q(n4914), .QN(n1102)
         );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n4670), .CK(CLK), .Q(n4913), .QN(n1103)
         );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n4671), .CK(CLK), .Q(n4912), .QN(n1104)
         );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n4672), .CK(CLK), .Q(n4911), .QN(n1105)
         );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n4673), .CK(CLK), .Q(n4910), .QN(n1106)
         );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n4674), .CK(CLK), .Q(n4909), .QN(n1107)
         );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n4675), .CK(CLK), .Q(n4908), .QN(n1108)
         );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n4676), .CK(CLK), .Q(n4907), .QN(n1109)
         );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n4677), .CK(CLK), .Q(n4906), .QN(n1110)
         );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n4678), .CK(CLK), .Q(n4905), .QN(n1111)
         );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n4679), .CK(CLK), .Q(n4904), .QN(n1112)
         );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n4680), .CK(CLK), .Q(n4903), .QN(n1113)
         );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n4681), .CK(CLK), .Q(n4902), .QN(n1114)
         );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n4682), .CK(CLK), .Q(n4901), .QN(n1115)
         );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n4683), .CK(CLK), .Q(n4900), .QN(n1116)
         );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n4684), .CK(CLK), .Q(n4899), .QN(n1117)
         );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n4685), .CK(CLK), .Q(n4898), .QN(n1118)
         );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n4686), .CK(CLK), .Q(n4897), .QN(n1119)
         );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n4687), .CK(CLK), .Q(n4896), .QN(n1120)
         );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n4688), .CK(CLK), .Q(n4895), .QN(n1121)
         );
  DFF_X1 \REGISTERS_reg[15][63]  ( .D(n4689), .CK(CLK), .Q(n5556), .QN(n1122)
         );
  DFF_X1 \REGISTERS_reg[15][62]  ( .D(n4690), .CK(CLK), .Q(n5555), .QN(n1123)
         );
  DFF_X1 \REGISTERS_reg[15][61]  ( .D(n4691), .CK(CLK), .Q(n5554), .QN(n1124)
         );
  DFF_X1 \REGISTERS_reg[15][60]  ( .D(n4692), .CK(CLK), .Q(n5553), .QN(n1125)
         );
  DFF_X1 \REGISTERS_reg[15][59]  ( .D(n4693), .CK(CLK), .Q(n5552), .QN(n1126)
         );
  DFF_X1 \REGISTERS_reg[15][58]  ( .D(n4694), .CK(CLK), .Q(n5551), .QN(n1127)
         );
  DFF_X1 \REGISTERS_reg[15][57]  ( .D(n4695), .CK(CLK), .Q(n5550), .QN(n1128)
         );
  DFF_X1 \REGISTERS_reg[15][56]  ( .D(n4696), .CK(CLK), .Q(n5549), .QN(n1129)
         );
  DFF_X1 \REGISTERS_reg[15][55]  ( .D(n4697), .CK(CLK), .Q(n5548), .QN(n1130)
         );
  DFF_X1 \REGISTERS_reg[15][54]  ( .D(n4698), .CK(CLK), .Q(n5547), .QN(n1131)
         );
  DFF_X1 \REGISTERS_reg[15][53]  ( .D(n4699), .CK(CLK), .Q(n5546), .QN(n1132)
         );
  DFF_X1 \REGISTERS_reg[15][52]  ( .D(n4700), .CK(CLK), .Q(n5545), .QN(n1133)
         );
  DFF_X1 \REGISTERS_reg[15][51]  ( .D(n4701), .CK(CLK), .Q(n5544), .QN(n1134)
         );
  DFF_X1 \REGISTERS_reg[15][50]  ( .D(n4702), .CK(CLK), .Q(n5543), .QN(n1135)
         );
  DFF_X1 \REGISTERS_reg[15][49]  ( .D(n4703), .CK(CLK), .Q(n5542), .QN(n1136)
         );
  DFF_X1 \REGISTERS_reg[15][48]  ( .D(n4704), .CK(CLK), .Q(n5541), .QN(n1137)
         );
  DFF_X1 \REGISTERS_reg[15][47]  ( .D(n4705), .CK(CLK), .Q(n5540), .QN(n1138)
         );
  DFF_X1 \REGISTERS_reg[15][46]  ( .D(n4706), .CK(CLK), .Q(n5539), .QN(n1139)
         );
  DFF_X1 \REGISTERS_reg[15][45]  ( .D(n4707), .CK(CLK), .Q(n5538), .QN(n1140)
         );
  DFF_X1 \REGISTERS_reg[15][44]  ( .D(n4708), .CK(CLK), .Q(n5537), .QN(n1141)
         );
  DFF_X1 \REGISTERS_reg[15][43]  ( .D(n4709), .CK(CLK), .Q(n5536), .QN(n1142)
         );
  DFF_X1 \REGISTERS_reg[15][42]  ( .D(n4710), .CK(CLK), .Q(n5535), .QN(n1143)
         );
  DFF_X1 \REGISTERS_reg[15][41]  ( .D(n4711), .CK(CLK), .Q(n5534), .QN(n1144)
         );
  DFF_X1 \REGISTERS_reg[15][40]  ( .D(n4712), .CK(CLK), .Q(n5533), .QN(n1145)
         );
  DFF_X1 \REGISTERS_reg[15][39]  ( .D(n4713), .CK(CLK), .Q(n5532), .QN(n1146)
         );
  DFF_X1 \REGISTERS_reg[15][38]  ( .D(n4714), .CK(CLK), .Q(n5531), .QN(n1147)
         );
  DFF_X1 \REGISTERS_reg[15][37]  ( .D(n4715), .CK(CLK), .Q(n5530), .QN(n1148)
         );
  DFF_X1 \REGISTERS_reg[15][36]  ( .D(n4716), .CK(CLK), .Q(n5529), .QN(n1149)
         );
  DFF_X1 \REGISTERS_reg[15][35]  ( .D(n4717), .CK(CLK), .Q(n5528), .QN(n1150)
         );
  DFF_X1 \REGISTERS_reg[15][34]  ( .D(n4718), .CK(CLK), .Q(n5527), .QN(n1151)
         );
  DFF_X1 \REGISTERS_reg[15][33]  ( .D(n4719), .CK(CLK), .Q(n5526), .QN(n1152)
         );
  DFF_X1 \REGISTERS_reg[15][32]  ( .D(n4720), .CK(CLK), .Q(n5525), .QN(n1153)
         );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n4721), .CK(CLK), .Q(n5524), .QN(n1154)
         );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n4722), .CK(CLK), .Q(n5523), .QN(n1155)
         );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n4723), .CK(CLK), .Q(n5522), .QN(n1156)
         );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n4724), .CK(CLK), .Q(n5521), .QN(n1157)
         );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n4725), .CK(CLK), .Q(n5520), .QN(n1158)
         );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n4726), .CK(CLK), .Q(n5519), .QN(n1159)
         );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n4727), .CK(CLK), .Q(n5518), .QN(n1160)
         );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n4728), .CK(CLK), .Q(n5517), .QN(n1161)
         );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n4729), .CK(CLK), .Q(n5516), .QN(n1162)
         );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n4730), .CK(CLK), .Q(n5515), .QN(n1163)
         );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n4731), .CK(CLK), .Q(n5514), .QN(n1164)
         );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n4732), .CK(CLK), .Q(n5513), .QN(n1165)
         );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n4733), .CK(CLK), .Q(n5512), .QN(n1166)
         );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n4734), .CK(CLK), .Q(n5511), .QN(n1167)
         );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n4735), .CK(CLK), .Q(n5510), .QN(n1168)
         );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n4736), .CK(CLK), .Q(n5509), .QN(n1169)
         );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n4737), .CK(CLK), .Q(n5508), .QN(n1170)
         );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n4738), .CK(CLK), .Q(n5507), .QN(n1171)
         );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n4739), .CK(CLK), .Q(n5506), .QN(n1172)
         );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n4740), .CK(CLK), .Q(n5505), .QN(n1173)
         );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n4741), .CK(CLK), .Q(n5504), .QN(n1174)
         );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n4742), .CK(CLK), .Q(n5503), .QN(n1175)
         );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n4743), .CK(CLK), .Q(n5502), .QN(n1176)
         );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n4744), .CK(CLK), .Q(n5501), .QN(n1177)
         );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n4745), .CK(CLK), .Q(n5500), .QN(n1178)
         );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n4746), .CK(CLK), .Q(n5499), .QN(n1179)
         );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n4747), .CK(CLK), .Q(n5498), .QN(n1180)
         );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n4748), .CK(CLK), .Q(n5497), .QN(n1181)
         );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n4749), .CK(CLK), .Q(n5496), .QN(n1182)
         );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n4750), .CK(CLK), .Q(n5495), .QN(n1183)
         );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n4751), .CK(CLK), .Q(n5494), .QN(n1184)
         );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n4752), .CK(CLK), .Q(n5493), .QN(n1185)
         );
  DFF_X1 \REGISTERS_reg[16][63]  ( .D(n4753), .CK(CLK), .Q(n8245), .QN(n5089)
         );
  DFF_X1 \OUT2_reg[63]  ( .D(n3601), .CK(CLK), .Q(OUT2[63]) );
  DFF_X1 \BUSOUT_reg[63]  ( .D(n8311), .CK(CLK), .Q(BUSOUT[63]), .QN(n7861) );
  DFF_X1 \REGISTERS_reg[16][62]  ( .D(n4754), .CK(CLK), .Q(n8246), .QN(n5088)
         );
  DFF_X1 \OUT2_reg[62]  ( .D(n3602), .CK(CLK), .Q(OUT2[62]) );
  DFF_X1 \BUSOUT_reg[62]  ( .D(n8312), .CK(CLK), .Q(BUSOUT[62]), .QN(n7862) );
  DFF_X1 \REGISTERS_reg[16][61]  ( .D(n4755), .CK(CLK), .Q(n8247), .QN(n5087)
         );
  DFF_X1 \OUT2_reg[61]  ( .D(n3603), .CK(CLK), .Q(OUT2[61]) );
  DFF_X1 \BUSOUT_reg[61]  ( .D(n8313), .CK(CLK), .Q(BUSOUT[61]), .QN(n7863) );
  DFF_X1 \REGISTERS_reg[16][60]  ( .D(n4756), .CK(CLK), .Q(n8248), .QN(n5086)
         );
  DFF_X1 \OUT2_reg[60]  ( .D(n3604), .CK(CLK), .Q(OUT2[60]) );
  DFF_X1 \BUSOUT_reg[60]  ( .D(n8314), .CK(CLK), .Q(BUSOUT[60]), .QN(n7864) );
  DFF_X1 \REGISTERS_reg[16][59]  ( .D(n4757), .CK(CLK), .Q(n8249), .QN(n5085)
         );
  DFF_X1 \OUT2_reg[59]  ( .D(n3605), .CK(CLK), .Q(OUT2[59]) );
  DFF_X1 \BUSOUT_reg[59]  ( .D(n8315), .CK(CLK), .Q(BUSOUT[59]), .QN(n7865) );
  DFF_X1 \REGISTERS_reg[16][58]  ( .D(n4758), .CK(CLK), .Q(n8250), .QN(n5084)
         );
  DFF_X1 \OUT2_reg[58]  ( .D(n3606), .CK(CLK), .Q(OUT2[58]) );
  DFF_X1 \BUSOUT_reg[58]  ( .D(n8316), .CK(CLK), .Q(BUSOUT[58]), .QN(n7866) );
  DFF_X1 \REGISTERS_reg[16][57]  ( .D(n4759), .CK(CLK), .Q(n8251), .QN(n5083)
         );
  DFF_X1 \OUT2_reg[57]  ( .D(n3607), .CK(CLK), .Q(OUT2[57]) );
  DFF_X1 \BUSOUT_reg[57]  ( .D(n8317), .CK(CLK), .Q(BUSOUT[57]), .QN(n7867) );
  DFF_X1 \REGISTERS_reg[16][56]  ( .D(n4760), .CK(CLK), .Q(n8252), .QN(n5082)
         );
  DFF_X1 \OUT2_reg[56]  ( .D(n3608), .CK(CLK), .Q(OUT2[56]) );
  DFF_X1 \BUSOUT_reg[56]  ( .D(n8318), .CK(CLK), .Q(BUSOUT[56]), .QN(n7868) );
  DFF_X1 \REGISTERS_reg[16][55]  ( .D(n4761), .CK(CLK), .Q(n8253), .QN(n5081)
         );
  DFF_X1 \OUT2_reg[55]  ( .D(n3609), .CK(CLK), .Q(OUT2[55]) );
  DFF_X1 \BUSOUT_reg[55]  ( .D(n8319), .CK(CLK), .Q(BUSOUT[55]), .QN(n7869) );
  DFF_X1 \REGISTERS_reg[16][54]  ( .D(n4762), .CK(CLK), .Q(n8254), .QN(n5080)
         );
  DFF_X1 \OUT2_reg[54]  ( .D(n3610), .CK(CLK), .Q(OUT2[54]) );
  DFF_X1 \BUSOUT_reg[54]  ( .D(n8320), .CK(CLK), .Q(BUSOUT[54]), .QN(n7870) );
  DFF_X1 \REGISTERS_reg[16][53]  ( .D(n4763), .CK(CLK), .Q(n8255), .QN(n5079)
         );
  DFF_X1 \OUT2_reg[53]  ( .D(n3611), .CK(CLK), .Q(OUT2[53]) );
  DFF_X1 \BUSOUT_reg[53]  ( .D(n8321), .CK(CLK), .Q(BUSOUT[53]), .QN(n7871) );
  DFF_X1 \REGISTERS_reg[16][52]  ( .D(n4764), .CK(CLK), .Q(n8256), .QN(n5078)
         );
  DFF_X1 \OUT2_reg[52]  ( .D(n3612), .CK(CLK), .Q(OUT2[52]) );
  DFF_X1 \BUSOUT_reg[52]  ( .D(n8322), .CK(CLK), .Q(BUSOUT[52]), .QN(n7872) );
  DFF_X1 \REGISTERS_reg[16][51]  ( .D(n4765), .CK(CLK), .Q(n8257), .QN(n5077)
         );
  DFF_X1 \OUT2_reg[51]  ( .D(n3613), .CK(CLK), .Q(OUT2[51]) );
  DFF_X1 \BUSOUT_reg[51]  ( .D(n8323), .CK(CLK), .Q(BUSOUT[51]), .QN(n7873) );
  DFF_X1 \REGISTERS_reg[16][50]  ( .D(n4766), .CK(CLK), .Q(n8258), .QN(n5076)
         );
  DFF_X1 \OUT2_reg[50]  ( .D(n3614), .CK(CLK), .Q(OUT2[50]) );
  DFF_X1 \BUSOUT_reg[50]  ( .D(n8324), .CK(CLK), .Q(BUSOUT[50]), .QN(n7874) );
  DFF_X1 \REGISTERS_reg[16][49]  ( .D(n4767), .CK(CLK), .Q(n8259), .QN(n5075)
         );
  DFF_X1 \OUT2_reg[49]  ( .D(n3615), .CK(CLK), .Q(OUT2[49]) );
  DFF_X1 \BUSOUT_reg[49]  ( .D(n8325), .CK(CLK), .Q(BUSOUT[49]), .QN(n7875) );
  DFF_X1 \REGISTERS_reg[16][48]  ( .D(n4768), .CK(CLK), .Q(n8260), .QN(n5074)
         );
  DFF_X1 \OUT2_reg[48]  ( .D(n3616), .CK(CLK), .Q(OUT2[48]) );
  DFF_X1 \BUSOUT_reg[48]  ( .D(n8326), .CK(CLK), .Q(BUSOUT[48]), .QN(n7876) );
  DFF_X1 \REGISTERS_reg[16][47]  ( .D(n4769), .CK(CLK), .Q(n8261), .QN(n5073)
         );
  DFF_X1 \OUT2_reg[47]  ( .D(n3617), .CK(CLK), .Q(OUT2[47]) );
  DFF_X1 \BUSOUT_reg[47]  ( .D(n8327), .CK(CLK), .Q(BUSOUT[47]), .QN(n7877) );
  DFF_X1 \REGISTERS_reg[16][46]  ( .D(n4770), .CK(CLK), .Q(n8262), .QN(n5072)
         );
  DFF_X1 \OUT2_reg[46]  ( .D(n3618), .CK(CLK), .Q(OUT2[46]) );
  DFF_X1 \BUSOUT_reg[46]  ( .D(n8328), .CK(CLK), .Q(BUSOUT[46]), .QN(n7878) );
  DFF_X1 \REGISTERS_reg[16][45]  ( .D(n4771), .CK(CLK), .Q(n8263), .QN(n5071)
         );
  DFF_X1 \OUT2_reg[45]  ( .D(n3619), .CK(CLK), .Q(OUT2[45]) );
  DFF_X1 \BUSOUT_reg[45]  ( .D(n8329), .CK(CLK), .Q(BUSOUT[45]), .QN(n7879) );
  DFF_X1 \REGISTERS_reg[16][44]  ( .D(n4772), .CK(CLK), .Q(n8264), .QN(n5070)
         );
  DFF_X1 \OUT2_reg[44]  ( .D(n3620), .CK(CLK), .Q(OUT2[44]) );
  DFF_X1 \BUSOUT_reg[44]  ( .D(n8330), .CK(CLK), .Q(BUSOUT[44]), .QN(n7880) );
  DFF_X1 \REGISTERS_reg[16][43]  ( .D(n4773), .CK(CLK), .Q(n8265), .QN(n5069)
         );
  DFF_X1 \OUT2_reg[43]  ( .D(n3621), .CK(CLK), .Q(OUT2[43]) );
  DFF_X1 \BUSOUT_reg[43]  ( .D(n8331), .CK(CLK), .Q(BUSOUT[43]), .QN(n7881) );
  DFF_X1 \REGISTERS_reg[16][42]  ( .D(n4774), .CK(CLK), .Q(n8266), .QN(n5068)
         );
  DFF_X1 \OUT2_reg[42]  ( .D(n3622), .CK(CLK), .Q(OUT2[42]) );
  DFF_X1 \BUSOUT_reg[42]  ( .D(n8332), .CK(CLK), .Q(BUSOUT[42]), .QN(n7882) );
  DFF_X1 \REGISTERS_reg[16][41]  ( .D(n4775), .CK(CLK), .Q(n8267), .QN(n5067)
         );
  DFF_X1 \OUT2_reg[41]  ( .D(n3623), .CK(CLK), .Q(OUT2[41]) );
  DFF_X1 \BUSOUT_reg[41]  ( .D(n8333), .CK(CLK), .Q(BUSOUT[41]), .QN(n7883) );
  DFF_X1 \REGISTERS_reg[16][40]  ( .D(n4776), .CK(CLK), .Q(n8268), .QN(n5066)
         );
  DFF_X1 \OUT2_reg[40]  ( .D(n3624), .CK(CLK), .Q(OUT2[40]) );
  DFF_X1 \BUSOUT_reg[40]  ( .D(n8334), .CK(CLK), .Q(BUSOUT[40]), .QN(n7884) );
  DFF_X1 \REGISTERS_reg[16][39]  ( .D(n4777), .CK(CLK), .Q(n8269), .QN(n5065)
         );
  DFF_X1 \OUT2_reg[39]  ( .D(n3625), .CK(CLK), .Q(OUT2[39]) );
  DFF_X1 \BUSOUT_reg[39]  ( .D(n8335), .CK(CLK), .Q(BUSOUT[39]), .QN(n7885) );
  DFF_X1 \REGISTERS_reg[16][38]  ( .D(n4778), .CK(CLK), .Q(n8270), .QN(n5064)
         );
  DFF_X1 \OUT2_reg[38]  ( .D(n3626), .CK(CLK), .Q(OUT2[38]) );
  DFF_X1 \BUSOUT_reg[38]  ( .D(n8336), .CK(CLK), .Q(BUSOUT[38]), .QN(n7886) );
  DFF_X1 \REGISTERS_reg[16][37]  ( .D(n4779), .CK(CLK), .Q(n8271), .QN(n5063)
         );
  DFF_X1 \OUT2_reg[37]  ( .D(n3627), .CK(CLK), .Q(OUT2[37]) );
  DFF_X1 \BUSOUT_reg[37]  ( .D(n8337), .CK(CLK), .Q(BUSOUT[37]), .QN(n7887) );
  DFF_X1 \REGISTERS_reg[16][36]  ( .D(n4780), .CK(CLK), .Q(n8272), .QN(n5062)
         );
  DFF_X1 \OUT2_reg[36]  ( .D(n3628), .CK(CLK), .Q(OUT2[36]) );
  DFF_X1 \BUSOUT_reg[36]  ( .D(n8338), .CK(CLK), .Q(BUSOUT[36]), .QN(n7888) );
  DFF_X1 \REGISTERS_reg[16][35]  ( .D(n4781), .CK(CLK), .Q(n8273), .QN(n5061)
         );
  DFF_X1 \OUT2_reg[35]  ( .D(n3629), .CK(CLK), .Q(OUT2[35]) );
  DFF_X1 \BUSOUT_reg[35]  ( .D(n8339), .CK(CLK), .Q(BUSOUT[35]), .QN(n7889) );
  DFF_X1 \REGISTERS_reg[16][34]  ( .D(n4782), .CK(CLK), .Q(n8274), .QN(n5060)
         );
  DFF_X1 \OUT2_reg[34]  ( .D(n3630), .CK(CLK), .Q(OUT2[34]) );
  DFF_X1 \BUSOUT_reg[34]  ( .D(n8340), .CK(CLK), .Q(BUSOUT[34]), .QN(n7890) );
  DFF_X1 \REGISTERS_reg[16][33]  ( .D(n4783), .CK(CLK), .Q(n8275), .QN(n5059)
         );
  DFF_X1 \OUT2_reg[33]  ( .D(n3631), .CK(CLK), .Q(OUT2[33]) );
  DFF_X1 \BUSOUT_reg[33]  ( .D(n8341), .CK(CLK), .Q(BUSOUT[33]), .QN(n7891) );
  DFF_X1 \REGISTERS_reg[16][32]  ( .D(n4784), .CK(CLK), .Q(n8276), .QN(n5058)
         );
  DFF_X1 \OUT2_reg[32]  ( .D(n3632), .CK(CLK), .Q(OUT2[32]) );
  DFF_X1 \BUSOUT_reg[32]  ( .D(n8342), .CK(CLK), .Q(BUSOUT[32]), .QN(n7892) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n4785), .CK(CLK), .Q(n8277), .QN(n5057)
         );
  DFF_X1 \OUT2_reg[31]  ( .D(n3633), .CK(CLK), .Q(OUT2[31]) );
  DFF_X1 \BUSOUT_reg[31]  ( .D(n8343), .CK(CLK), .Q(BUSOUT[31]), .QN(n7893) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n4786), .CK(CLK), .Q(n8278), .QN(n5056)
         );
  DFF_X1 \OUT2_reg[30]  ( .D(n3634), .CK(CLK), .Q(OUT2[30]) );
  DFF_X1 \BUSOUT_reg[30]  ( .D(n8344), .CK(CLK), .Q(BUSOUT[30]), .QN(n7894) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n4787), .CK(CLK), .Q(n8279), .QN(n5055)
         );
  DFF_X1 \OUT2_reg[29]  ( .D(n3635), .CK(CLK), .Q(OUT2[29]) );
  DFF_X1 \BUSOUT_reg[29]  ( .D(n8345), .CK(CLK), .Q(BUSOUT[29]), .QN(n7895) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n4788), .CK(CLK), .Q(n8280), .QN(n5054)
         );
  DFF_X1 \OUT2_reg[28]  ( .D(n3636), .CK(CLK), .Q(OUT2[28]) );
  DFF_X1 \BUSOUT_reg[28]  ( .D(n8346), .CK(CLK), .Q(BUSOUT[28]), .QN(n7896) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n4789), .CK(CLK), .Q(n8281), .QN(n5053)
         );
  DFF_X1 \OUT2_reg[27]  ( .D(n3637), .CK(CLK), .Q(OUT2[27]) );
  DFF_X1 \BUSOUT_reg[27]  ( .D(n8347), .CK(CLK), .Q(BUSOUT[27]), .QN(n7897) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n4790), .CK(CLK), .Q(n8282), .QN(n5052)
         );
  DFF_X1 \OUT2_reg[26]  ( .D(n3638), .CK(CLK), .Q(OUT2[26]) );
  DFF_X1 \BUSOUT_reg[26]  ( .D(n8348), .CK(CLK), .Q(BUSOUT[26]), .QN(n7898) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n4791), .CK(CLK), .Q(n8283), .QN(n5051)
         );
  DFF_X1 \OUT2_reg[25]  ( .D(n3639), .CK(CLK), .Q(OUT2[25]) );
  DFF_X1 \BUSOUT_reg[25]  ( .D(n8349), .CK(CLK), .Q(BUSOUT[25]), .QN(n7899) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n4792), .CK(CLK), .Q(n8284), .QN(n5050)
         );
  DFF_X1 \OUT2_reg[24]  ( .D(n3640), .CK(CLK), .Q(OUT2[24]) );
  DFF_X1 \BUSOUT_reg[24]  ( .D(n8350), .CK(CLK), .Q(BUSOUT[24]), .QN(n7900) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n4793), .CK(CLK), .Q(n8285), .QN(n5049)
         );
  DFF_X1 \OUT2_reg[23]  ( .D(n3641), .CK(CLK), .Q(OUT2[23]) );
  DFF_X1 \BUSOUT_reg[23]  ( .D(n8351), .CK(CLK), .Q(BUSOUT[23]), .QN(n7901) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n4794), .CK(CLK), .Q(n8286), .QN(n5048)
         );
  DFF_X1 \OUT2_reg[22]  ( .D(n3642), .CK(CLK), .Q(OUT2[22]) );
  DFF_X1 \BUSOUT_reg[22]  ( .D(n8352), .CK(CLK), .Q(BUSOUT[22]), .QN(n7902) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n4795), .CK(CLK), .Q(n8287), .QN(n5047)
         );
  DFF_X1 \OUT2_reg[21]  ( .D(n3643), .CK(CLK), .Q(OUT2[21]) );
  DFF_X1 \BUSOUT_reg[21]  ( .D(n8353), .CK(CLK), .Q(BUSOUT[21]), .QN(n7903) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n4796), .CK(CLK), .Q(n8288), .QN(n5046)
         );
  DFF_X1 \OUT2_reg[20]  ( .D(n3644), .CK(CLK), .Q(OUT2[20]) );
  DFF_X1 \BUSOUT_reg[20]  ( .D(n8354), .CK(CLK), .Q(BUSOUT[20]), .QN(n7904) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n4797), .CK(CLK), .Q(n8289), .QN(n5045)
         );
  DFF_X1 \OUT2_reg[19]  ( .D(n3645), .CK(CLK), .Q(OUT2[19]) );
  DFF_X1 \BUSOUT_reg[19]  ( .D(n8355), .CK(CLK), .Q(BUSOUT[19]), .QN(n7905) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n4798), .CK(CLK), .Q(n8290), .QN(n5044)
         );
  DFF_X1 \OUT2_reg[18]  ( .D(n3646), .CK(CLK), .Q(OUT2[18]) );
  DFF_X1 \BUSOUT_reg[18]  ( .D(n8356), .CK(CLK), .Q(BUSOUT[18]), .QN(n7906) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n4799), .CK(CLK), .Q(n8291), .QN(n5043)
         );
  DFF_X1 \OUT2_reg[17]  ( .D(n3647), .CK(CLK), .Q(OUT2[17]) );
  DFF_X1 \BUSOUT_reg[17]  ( .D(n8357), .CK(CLK), .Q(BUSOUT[17]), .QN(n7907) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n4800), .CK(CLK), .Q(n8292), .QN(n5042)
         );
  DFF_X1 \OUT2_reg[16]  ( .D(n3648), .CK(CLK), .Q(OUT2[16]) );
  DFF_X1 \BUSOUT_reg[16]  ( .D(n8358), .CK(CLK), .Q(BUSOUT[16]), .QN(n7908) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n4801), .CK(CLK), .Q(n8293), .QN(n5041)
         );
  DFF_X1 \OUT2_reg[15]  ( .D(n3649), .CK(CLK), .Q(OUT2[15]) );
  DFF_X1 \BUSOUT_reg[15]  ( .D(n8359), .CK(CLK), .Q(BUSOUT[15]), .QN(n7909) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n4802), .CK(CLK), .Q(n8294), .QN(n5040)
         );
  DFF_X1 \OUT2_reg[14]  ( .D(n3650), .CK(CLK), .Q(OUT2[14]) );
  DFF_X1 \BUSOUT_reg[14]  ( .D(n8360), .CK(CLK), .Q(BUSOUT[14]), .QN(n7910) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n4803), .CK(CLK), .Q(n8295), .QN(n5039)
         );
  DFF_X1 \OUT2_reg[13]  ( .D(n3651), .CK(CLK), .Q(OUT2[13]) );
  DFF_X1 \BUSOUT_reg[13]  ( .D(n8361), .CK(CLK), .Q(BUSOUT[13]), .QN(n7911) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n4804), .CK(CLK), .Q(n8296), .QN(n5038)
         );
  DFF_X1 \OUT2_reg[12]  ( .D(n3652), .CK(CLK), .Q(OUT2[12]) );
  DFF_X1 \BUSOUT_reg[12]  ( .D(n8362), .CK(CLK), .Q(BUSOUT[12]), .QN(n7912) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n4805), .CK(CLK), .Q(n8297), .QN(n5037)
         );
  DFF_X1 \OUT2_reg[11]  ( .D(n3653), .CK(CLK), .Q(OUT2[11]) );
  DFF_X1 \BUSOUT_reg[11]  ( .D(n8363), .CK(CLK), .Q(BUSOUT[11]), .QN(n7913) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n4806), .CK(CLK), .Q(n8298), .QN(n5036)
         );
  DFF_X1 \OUT2_reg[10]  ( .D(n3654), .CK(CLK), .Q(OUT2[10]) );
  DFF_X1 \BUSOUT_reg[10]  ( .D(n8364), .CK(CLK), .Q(BUSOUT[10]), .QN(n7914) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n4807), .CK(CLK), .Q(n8299), .QN(n5035)
         );
  DFF_X1 \OUT2_reg[9]  ( .D(n3655), .CK(CLK), .Q(OUT2[9]) );
  DFF_X1 \BUSOUT_reg[9]  ( .D(n8365), .CK(CLK), .Q(BUSOUT[9]), .QN(n7915) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n4808), .CK(CLK), .Q(n8300), .QN(n5034)
         );
  DFF_X1 \OUT2_reg[8]  ( .D(n3656), .CK(CLK), .Q(OUT2[8]) );
  DFF_X1 \BUSOUT_reg[8]  ( .D(n8366), .CK(CLK), .Q(BUSOUT[8]), .QN(n7916) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n4809), .CK(CLK), .Q(n8301), .QN(n5033)
         );
  DFF_X1 \OUT2_reg[7]  ( .D(n3657), .CK(CLK), .Q(OUT2[7]) );
  DFF_X1 \BUSOUT_reg[7]  ( .D(n8367), .CK(CLK), .Q(BUSOUT[7]), .QN(n7917) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n4810), .CK(CLK), .Q(n8302), .QN(n5032)
         );
  DFF_X1 \OUT2_reg[6]  ( .D(n3658), .CK(CLK), .Q(OUT2[6]) );
  DFF_X1 \BUSOUT_reg[6]  ( .D(n8368), .CK(CLK), .Q(BUSOUT[6]), .QN(n7918) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n4811), .CK(CLK), .Q(n8303), .QN(n5031)
         );
  DFF_X1 \OUT2_reg[5]  ( .D(n3659), .CK(CLK), .Q(OUT2[5]) );
  DFF_X1 \BUSOUT_reg[5]  ( .D(n8369), .CK(CLK), .Q(BUSOUT[5]), .QN(n7919) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n4812), .CK(CLK), .Q(n8304), .QN(n5030)
         );
  DFF_X1 \OUT2_reg[4]  ( .D(n3660), .CK(CLK), .Q(OUT2[4]) );
  DFF_X1 \BUSOUT_reg[4]  ( .D(n8370), .CK(CLK), .Q(BUSOUT[4]), .QN(n7920) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n4813), .CK(CLK), .Q(n8305), .QN(n5029)
         );
  DFF_X1 \OUT2_reg[3]  ( .D(n3661), .CK(CLK), .Q(OUT2[3]) );
  DFF_X1 \BUSOUT_reg[3]  ( .D(n8371), .CK(CLK), .Q(BUSOUT[3]), .QN(n7921) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n4814), .CK(CLK), .Q(n8306), .QN(n5028)
         );
  DFF_X1 \OUT2_reg[2]  ( .D(n3662), .CK(CLK), .Q(OUT2[2]) );
  DFF_X1 \BUSOUT_reg[2]  ( .D(n8372), .CK(CLK), .Q(BUSOUT[2]), .QN(n7922) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n4815), .CK(CLK), .Q(n8307), .QN(n5027)
         );
  DFF_X1 \OUT2_reg[1]  ( .D(n3663), .CK(CLK), .Q(OUT2[1]) );
  DFF_X1 \BUSOUT_reg[1]  ( .D(n8373), .CK(CLK), .Q(BUSOUT[1]), .QN(n7923) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n4816), .CK(CLK), .Q(n8308), .QN(n5026)
         );
  DFF_X1 \OUT2_reg[0]  ( .D(n3664), .CK(CLK), .Q(OUT2[0]) );
  DFF_X1 \BUSOUT_reg[0]  ( .D(n8374), .CK(CLK), .Q(BUSOUT[0]), .QN(n7924) );
  DFF_X1 \OUT1_reg[63]  ( .D(n3665), .CK(CLK), .Q(OUT1[63]) );
  DFF_X1 \OUT1_reg[62]  ( .D(n3666), .CK(CLK), .Q(OUT1[62]) );
  DFF_X1 \OUT1_reg[61]  ( .D(n3667), .CK(CLK), .Q(OUT1[61]) );
  DFF_X1 \OUT1_reg[60]  ( .D(n3668), .CK(CLK), .Q(OUT1[60]) );
  DFF_X1 \OUT1_reg[59]  ( .D(n3669), .CK(CLK), .Q(OUT1[59]) );
  DFF_X1 \OUT1_reg[58]  ( .D(n3670), .CK(CLK), .Q(OUT1[58]) );
  DFF_X1 \OUT1_reg[57]  ( .D(n3671), .CK(CLK), .Q(OUT1[57]) );
  DFF_X1 \OUT1_reg[56]  ( .D(n3672), .CK(CLK), .Q(OUT1[56]) );
  DFF_X1 \OUT1_reg[55]  ( .D(n3673), .CK(CLK), .Q(OUT1[55]) );
  DFF_X1 \OUT1_reg[54]  ( .D(n3674), .CK(CLK), .Q(OUT1[54]) );
  DFF_X1 \OUT1_reg[53]  ( .D(n3675), .CK(CLK), .Q(OUT1[53]) );
  DFF_X1 \OUT1_reg[52]  ( .D(n3676), .CK(CLK), .Q(OUT1[52]) );
  DFF_X1 \OUT1_reg[51]  ( .D(n3677), .CK(CLK), .Q(OUT1[51]) );
  DFF_X1 \OUT1_reg[50]  ( .D(n3678), .CK(CLK), .Q(OUT1[50]) );
  DFF_X1 \OUT1_reg[49]  ( .D(n3679), .CK(CLK), .Q(OUT1[49]) );
  DFF_X1 \OUT1_reg[48]  ( .D(n3680), .CK(CLK), .Q(OUT1[48]) );
  DFF_X1 \OUT1_reg[47]  ( .D(n3681), .CK(CLK), .Q(OUT1[47]) );
  DFF_X1 \OUT1_reg[46]  ( .D(n3682), .CK(CLK), .Q(OUT1[46]) );
  DFF_X1 \OUT1_reg[45]  ( .D(n3683), .CK(CLK), .Q(OUT1[45]) );
  DFF_X1 \OUT1_reg[44]  ( .D(n3684), .CK(CLK), .Q(OUT1[44]) );
  DFF_X1 \OUT1_reg[43]  ( .D(n3685), .CK(CLK), .Q(OUT1[43]) );
  DFF_X1 \OUT1_reg[42]  ( .D(n3686), .CK(CLK), .Q(OUT1[42]) );
  DFF_X1 \OUT1_reg[41]  ( .D(n3687), .CK(CLK), .Q(OUT1[41]) );
  DFF_X1 \OUT1_reg[40]  ( .D(n3688), .CK(CLK), .Q(OUT1[40]) );
  DFF_X1 \OUT1_reg[39]  ( .D(n3689), .CK(CLK), .Q(OUT1[39]) );
  DFF_X1 \OUT1_reg[38]  ( .D(n3690), .CK(CLK), .Q(OUT1[38]) );
  DFF_X1 \OUT1_reg[37]  ( .D(n3691), .CK(CLK), .Q(OUT1[37]) );
  DFF_X1 \OUT1_reg[36]  ( .D(n3692), .CK(CLK), .Q(OUT1[36]) );
  DFF_X1 \OUT1_reg[35]  ( .D(n3693), .CK(CLK), .Q(OUT1[35]) );
  DFF_X1 \OUT1_reg[34]  ( .D(n3694), .CK(CLK), .Q(OUT1[34]) );
  DFF_X1 \OUT1_reg[33]  ( .D(n3695), .CK(CLK), .Q(OUT1[33]) );
  DFF_X1 \OUT1_reg[32]  ( .D(n3696), .CK(CLK), .Q(OUT1[32]) );
  DFF_X1 \OUT1_reg[31]  ( .D(n3697), .CK(CLK), .Q(OUT1[31]) );
  DFF_X1 \OUT1_reg[30]  ( .D(n3698), .CK(CLK), .Q(OUT1[30]) );
  DFF_X1 \OUT1_reg[29]  ( .D(n3699), .CK(CLK), .Q(OUT1[29]) );
  DFF_X1 \OUT1_reg[28]  ( .D(n3700), .CK(CLK), .Q(OUT1[28]) );
  DFF_X1 \OUT1_reg[27]  ( .D(n3701), .CK(CLK), .Q(OUT1[27]) );
  DFF_X1 \OUT1_reg[26]  ( .D(n3702), .CK(CLK), .Q(OUT1[26]) );
  DFF_X1 \OUT1_reg[25]  ( .D(n3703), .CK(CLK), .Q(OUT1[25]) );
  DFF_X1 \OUT1_reg[24]  ( .D(n3704), .CK(CLK), .Q(OUT1[24]) );
  DFF_X1 \OUT1_reg[23]  ( .D(n3705), .CK(CLK), .Q(OUT1[23]) );
  DFF_X1 \OUT1_reg[22]  ( .D(n3706), .CK(CLK), .Q(OUT1[22]) );
  DFF_X1 \OUT1_reg[21]  ( .D(n3707), .CK(CLK), .Q(OUT1[21]) );
  DFF_X1 \OUT1_reg[20]  ( .D(n3708), .CK(CLK), .Q(OUT1[20]) );
  DFF_X1 \OUT1_reg[19]  ( .D(n3709), .CK(CLK), .Q(OUT1[19]) );
  DFF_X1 \OUT1_reg[18]  ( .D(n3710), .CK(CLK), .Q(OUT1[18]) );
  DFF_X1 \OUT1_reg[17]  ( .D(n3711), .CK(CLK), .Q(OUT1[17]) );
  DFF_X1 \OUT1_reg[16]  ( .D(n3712), .CK(CLK), .Q(OUT1[16]) );
  DFF_X1 \OUT1_reg[15]  ( .D(n3713), .CK(CLK), .Q(OUT1[15]) );
  DFF_X1 \OUT1_reg[14]  ( .D(n3714), .CK(CLK), .Q(OUT1[14]) );
  DFF_X1 \OUT1_reg[13]  ( .D(n3715), .CK(CLK), .Q(OUT1[13]) );
  DFF_X1 \OUT1_reg[12]  ( .D(n3716), .CK(CLK), .Q(OUT1[12]) );
  DFF_X1 \OUT1_reg[11]  ( .D(n3717), .CK(CLK), .Q(OUT1[11]) );
  DFF_X1 \OUT1_reg[10]  ( .D(n3718), .CK(CLK), .Q(OUT1[10]) );
  DFF_X1 \OUT1_reg[9]  ( .D(n3719), .CK(CLK), .Q(OUT1[9]) );
  DFF_X1 \OUT1_reg[8]  ( .D(n3720), .CK(CLK), .Q(OUT1[8]) );
  DFF_X1 \OUT1_reg[7]  ( .D(n3721), .CK(CLK), .Q(OUT1[7]) );
  DFF_X1 \OUT1_reg[6]  ( .D(n3722), .CK(CLK), .Q(OUT1[6]) );
  DFF_X1 \OUT1_reg[5]  ( .D(n3723), .CK(CLK), .Q(OUT1[5]) );
  DFF_X1 \OUT1_reg[4]  ( .D(n3724), .CK(CLK), .Q(OUT1[4]) );
  DFF_X1 \OUT1_reg[3]  ( .D(n3725), .CK(CLK), .Q(OUT1[3]) );
  DFF_X1 \OUT1_reg[2]  ( .D(n3726), .CK(CLK), .Q(OUT1[2]) );
  DFF_X1 \OUT1_reg[1]  ( .D(n3727), .CK(CLK), .Q(OUT1[1]) );
  DFF_X1 \OUT1_reg[0]  ( .D(n3728), .CK(CLK), .Q(OUT1[0]) );
  FA_X1 \r631/U1_1  ( .A(SWP[1]), .B(n8310), .CI(\r631/carry[1] ), .CO(
        \r631/carry[2] ), .S(N924) );
  FA_X1 \r631/U1_2  ( .A(SWP[2]), .B(n8310), .CI(\r631/carry[2] ), .CO(
        \r631/carry[3] ), .S(N925) );
  FA_X1 \r631/U1_3  ( .A(SWP[3]), .B(\r631/carry[1] ), .CI(\r631/carry[3] ), 
        .CO(\r631/carry[4] ), .S(N926) );
  FA_X1 \r631/U1_4  ( .A(SWP[4]), .B(\r631/carry[1] ), .CI(\r631/carry[4] ), 
        .S(N927) );
  FA_X1 \r646/U1_1  ( .A(\U3/U199/Z_1 ), .B(\U3/U200/Z_1 ), .CI(n5854), .CO(
        \r646/carry[2] ), .S(N555) );
  FA_X1 \r646/U1_2  ( .A(\U3/U199/Z_2 ), .B(\U3/U200/Z_2 ), .CI(
        \r646/carry[2] ), .CO(\r646/carry[3] ), .S(N556) );
  FA_X1 \r646/U1_3  ( .A(\U3/U199/Z_3 ), .B(\U3/U200/Z_3 ), .CI(
        \r646/carry[3] ), .CO(\r646/carry[4] ), .S(N557) );
  FA_X1 \r642/U1_1  ( .A(\U3/U199/Z_1 ), .B(\U3/U200/Z_1 ), .CI(n5853), .CO(
        \r642/carry[2] ), .S(N332) );
  FA_X1 \r642/U1_2  ( .A(\U3/U199/Z_2 ), .B(\U3/U200/Z_2 ), .CI(
        \r642/carry[2] ), .CO(\r642/carry[3] ), .S(N333) );
  FA_X1 \r642/U1_3  ( .A(\U3/U199/Z_3 ), .B(\U3/U200/Z_3 ), .CI(
        \r642/carry[3] ), .CO(\r642/carry[4] ), .S(N334) );
  FA_X1 \r638/U1_1  ( .A(\U3/U195/Z_1 ), .B(\U3/U196/Z_1 ), .CI(n5558), .CO(
        \r638/carry[2] ), .S(N433) );
  FA_X1 \r638/U1_2  ( .A(\U3/U195/Z_2 ), .B(\U3/U196/Z_2 ), .CI(
        \r638/carry[2] ), .CO(\r638/carry[3] ), .S(N434) );
  FA_X1 \r638/U1_3  ( .A(\U3/U195/Z_3 ), .B(\U3/U196/Z_3 ), .CI(
        \r638/carry[3] ), .CO(\r638/carry[4] ), .S(N435) );
  FA_X1 \r507/U1_1  ( .A(\U3/U201/Z_1 ), .B(\U3/U202/Z_1 ), .CI(n5557), .CO(
        \r507/carry[2] ), .S(N208) );
  FA_X1 \r507/U1_2  ( .A(\U3/U201/Z_2 ), .B(\U3/U202/Z_2 ), .CI(
        \r507/carry[2] ), .CO(\r507/carry[3] ), .S(N209) );
  FA_X1 \r507/U1_3  ( .A(\U3/U201/Z_3 ), .B(\U3/U202/Z_3 ), .CI(
        \r507/carry[3] ), .CO(\r507/carry[4] ), .S(N210) );
  FA_X1 \r467/U1_1  ( .A(ADD_WR[1]), .B(CWP[1]), .CI(n5859), .CO(
        \r467/carry[2] ), .S(N560) );
  FA_X1 \r467/U1_2  ( .A(ADD_WR[2]), .B(CWP[2]), .CI(\r467/carry[2] ), .CO(
        \r467/carry[3] ), .S(N561) );
  FA_X1 \r467/U1_3  ( .A(ADD_WR[3]), .B(CWP[3]), .CI(\r467/carry[3] ), .CO(
        \r467/carry[4] ), .S(N562) );
  OR2_X1 U3676 ( .A1(FILL), .A2(RST), .ZN(n4959) );
  AND3_X1 U3677 ( .A1(n6467), .A2(n5877), .A3(n6461), .ZN(n4960) );
  AND3_X1 U3678 ( .A1(n7243), .A2(n7244), .A3(n7242), .ZN(n5218) );
  AND3_X1 U3679 ( .A1(n5851), .A2(n7244), .A3(n7251), .ZN(n5219) );
  AND3_X1 U3680 ( .A1(n7245), .A2(N333), .A3(n7254), .ZN(n5220) );
  AND3_X1 U3681 ( .A1(n7788), .A2(n7789), .A3(n7787), .ZN(n5221) );
  AND3_X1 U3682 ( .A1(n5852), .A2(n7789), .A3(n7797), .ZN(n5222) );
  AND3_X1 U3683 ( .A1(n7790), .A2(N434), .A3(n7800), .ZN(n5223) );
  AND2_X1 U3684 ( .A1(n6469), .A2(n6463), .ZN(n5224) );
  AND3_X1 U3685 ( .A1(n7245), .A2(N333), .A3(n7246), .ZN(n5225) );
  AND3_X1 U3686 ( .A1(n7790), .A2(N434), .A3(n7791), .ZN(n5226) );
  AND4_X1 U3687 ( .A1(n7254), .A2(n7248), .A3(n7247), .A4(n7257), .ZN(n5227)
         );
  AND4_X1 U3688 ( .A1(n7800), .A2(n7793), .A3(n7792), .A4(n7803), .ZN(n5228)
         );
  OR2_X1 U3689 ( .A1(RST), .A2(n1327), .ZN(n5229) );
  OR3_X1 U3690 ( .A1(n6738), .A2(RST), .A3(n7259), .ZN(n5230) );
  OR3_X1 U3691 ( .A1(n7283), .A2(RST), .A3(n7805), .ZN(n5231) );
  AND3_X1 U3692 ( .A1(n7242), .A2(n7243), .A3(N332), .ZN(n5232) );
  AND3_X1 U3693 ( .A1(n7245), .A2(n7247), .A3(n7254), .ZN(n5233) );
  AND3_X1 U3694 ( .A1(n7787), .A2(n7788), .A3(N433), .ZN(n5234) );
  AND3_X1 U3695 ( .A1(n7790), .A2(n7792), .A3(n7800), .ZN(n5235) );
  AND2_X1 U3696 ( .A1(\U3/U202/Z_0 ), .A2(\U3/U201/Z_0 ), .ZN(n5557) );
  AND2_X1 U3697 ( .A1(\U3/U196/Z_0 ), .A2(\U3/U195/Z_0 ), .ZN(n5558) );
  AND2_X4 U3698 ( .A1(n6465), .A2(n6471), .ZN(n5895) );
  AND2_X4 U3699 ( .A1(n6463), .A2(n6471), .ZN(n5894) );
  AND2_X4 U3700 ( .A1(n7249), .A2(n7248), .ZN(n6726) );
  AND2_X4 U3701 ( .A1(n7794), .A2(n7793), .ZN(n7271) );
  AND3_X4 U3702 ( .A1(n7790), .A2(n7792), .A3(n7791), .ZN(n7274) );
  AND3_X4 U3703 ( .A1(N433), .A2(n5852), .A3(n7797), .ZN(n7279) );
  AND3_X4 U3704 ( .A1(n7245), .A2(n7247), .A3(n7246), .ZN(n6729) );
  AND3_X4 U3705 ( .A1(N332), .A2(n5851), .A3(n7251), .ZN(n6734) );
  NAND2_X4 U3706 ( .A1(n7794), .A2(n7790), .ZN(n7278) );
  AND2_X4 U3707 ( .A1(n6461), .A2(n6462), .ZN(n5880) );
  NAND2_X4 U3708 ( .A1(n6467), .A2(n6471), .ZN(n5891) );
  NAND2_X4 U3709 ( .A1(n7249), .A2(n7245), .ZN(n6733) );
  NAND2_X4 U3710 ( .A1(n6466), .A2(n6462), .ZN(n5882) );
  NAND2_X4 U3711 ( .A1(n6469), .A2(n6462), .ZN(n5886) );
  INV_X4 U3712 ( .A(n5234), .ZN(n5815) );
  INV_X4 U3713 ( .A(n5235), .ZN(n5816) );
  INV_X4 U3714 ( .A(n5232), .ZN(n5817) );
  INV_X4 U3715 ( .A(n5233), .ZN(n5818) );
  NAND2_X4 U3716 ( .A1(n7797), .A2(n7791), .ZN(n7277) );
  NAND2_X4 U3717 ( .A1(n5864), .A2(n7788), .ZN(n7282) );
  NAND2_X4 U3718 ( .A1(n7251), .A2(n7246), .ZN(n6732) );
  NAND2_X4 U3719 ( .A1(n5856), .A2(n7243), .ZN(n6737) );
  AND2_X4 U3720 ( .A1(n6461), .A2(n6465), .ZN(n5885) );
  AND2_X4 U3721 ( .A1(n6466), .A2(n6465), .ZN(n5889) );
  INV_X4 U3722 ( .A(n5224), .ZN(n5819) );
  NAND2_X4 U3723 ( .A1(n6469), .A2(n6465), .ZN(n5890) );
  INV_X4 U3724 ( .A(n5226), .ZN(n5820) );
  NAND2_X4 U3725 ( .A1(n6466), .A2(n6463), .ZN(n5881) );
  INV_X4 U3726 ( .A(n5225), .ZN(n5821) );
  INV_X4 U3727 ( .A(n5860), .ZN(n5877) );
  AND2_X4 U3728 ( .A1(n7798), .A2(n7790), .ZN(n7275) );
  AND2_X4 U3729 ( .A1(n7800), .A2(n7797), .ZN(n7280) );
  AND2_X4 U3730 ( .A1(n7252), .A2(n7245), .ZN(n6730) );
  AND2_X4 U3731 ( .A1(n7254), .A2(n7251), .ZN(n6735) );
  AND3_X4 U3732 ( .A1(n7246), .A2(n7247), .A3(n7248), .ZN(n6727) );
  AND3_X4 U3733 ( .A1(n7791), .A2(n7792), .A3(n7793), .ZN(n7272) );
  NAND2_X4 U3734 ( .A1(n7252), .A2(n7248), .ZN(n6740) );
  NAND2_X4 U3735 ( .A1(n7798), .A2(n7793), .ZN(n7285) );
  AND2_X4 U3736 ( .A1(n6462), .A2(n6471), .ZN(n5893) );
  NAND2_X4 U3737 ( .A1(n5870), .A2(n6455), .ZN(n5872) );
  INV_X4 U3738 ( .A(n5220), .ZN(n5822) );
  INV_X4 U3739 ( .A(n5221), .ZN(n5823) );
  INV_X4 U3740 ( .A(n5222), .ZN(n5824) );
  INV_X4 U3741 ( .A(n5223), .ZN(n5825) );
  INV_X4 U3742 ( .A(n5227), .ZN(n5826) );
  INV_X4 U3743 ( .A(n5228), .ZN(n5827) );
  INV_X4 U3744 ( .A(n5218), .ZN(n5828) );
  INV_X4 U3745 ( .A(n5219), .ZN(n5829) );
  INV_X4 U3746 ( .A(n7804), .ZN(n7283) );
  AND2_X4 U3747 ( .A1(n6466), .A2(n6467), .ZN(n5884) );
  AND2_X4 U3748 ( .A1(n6467), .A2(n6469), .ZN(n5888) );
  AND2_X4 U3749 ( .A1(n6461), .A2(n6463), .ZN(n5879) );
  INV_X4 U3750 ( .A(n4960), .ZN(n5830) );
  AND3_X4 U3751 ( .A1(n6596), .A2(n6455), .A3(n6597), .ZN(n6532) );
  NAND2_X4 U3752 ( .A1(n1322), .A2(n6455), .ZN(n5870) );
  INV_X4 U3753 ( .A(n7258), .ZN(n6738) );
  INV_X4 U3754 ( .A(n4959), .ZN(n5831) );
  INV_X4 U3755 ( .A(n5230), .ZN(n5832) );
  INV_X4 U3756 ( .A(n5231), .ZN(n5833) );
  INV_X4 U3757 ( .A(n5229), .ZN(n5834) );
  INV_X1 U3758 ( .A(n6632), .ZN(n5835) );
  INV_X4 U3759 ( .A(n5835), .ZN(n5836) );
  INV_X1 U3760 ( .A(n6636), .ZN(n5837) );
  INV_X4 U3761 ( .A(n5837), .ZN(n5838) );
  INV_X1 U3762 ( .A(n6646), .ZN(n5839) );
  INV_X4 U3763 ( .A(n5839), .ZN(n5840) );
  INV_X1 U3764 ( .A(n6649), .ZN(n5841) );
  INV_X4 U3765 ( .A(n5841), .ZN(n5842) );
  INV_X1 U3766 ( .A(n6601), .ZN(n5843) );
  INV_X4 U3767 ( .A(n5843), .ZN(n5844) );
  INV_X1 U3768 ( .A(n6607), .ZN(n5845) );
  INV_X4 U3769 ( .A(n5845), .ZN(n5846) );
  INV_X1 U3770 ( .A(n6620), .ZN(n5847) );
  INV_X4 U3771 ( .A(n5847), .ZN(n5848) );
  INV_X1 U3772 ( .A(n6624), .ZN(n5849) );
  INV_X4 U3773 ( .A(n5849), .ZN(n5850) );
  AOI221_X4 U3774 ( .B1(n6627), .B2(n6635), .C1(n6463), .C2(n6653), .A(RST), 
        .ZN(n6652) );
  AOI221_X4 U3775 ( .B1(n4960), .B2(n6475), .C1(n6600), .C2(n6638), .A(RST), 
        .ZN(n6656) );
  AOI211_X4 U3776 ( .C1(n6467), .C2(n6613), .A(n6615), .B(RST), .ZN(n6614) );
  AOI211_X4 U3777 ( .C1(n6467), .C2(n6640), .A(n6642), .B(RST), .ZN(n6641) );
  AOI221_X4 U3778 ( .B1(n6605), .B2(n6612), .C1(n6463), .C2(n6613), .A(RST), 
        .ZN(n6611) );
  AOI221_X4 U3779 ( .B1(n6627), .B2(n6605), .C1(n6463), .C2(n6628), .A(RST), 
        .ZN(n6626) );
  AOI221_X4 U3780 ( .B1(n6600), .B2(n6609), .C1(n6467), .C2(n6628), .A(RST), 
        .ZN(n6630) );
  AOI221_X4 U3781 ( .B1(n6612), .B2(n6635), .C1(n6463), .C2(n6640), .A(RST), 
        .ZN(n6639) );
  INV_X1 U3782 ( .A(n5866), .ZN(N914) );
  XNOR2_X1 U3783 ( .A(n6629), .B(n5867), .ZN(n7263) );
  XNOR2_X1 U3784 ( .A(\U3/U200/Z_0 ), .B(\U3/U199/Z_0 ), .ZN(n5867) );
  XNOR2_X1 U3785 ( .A(n6598), .B(n5868), .ZN(n7265) );
  XNOR2_X1 U3786 ( .A(\U3/U200/Z_4 ), .B(\r646/carry[4] ), .ZN(n5868) );
  XOR2_X1 U3787 ( .A(\U3/U200/Z_0 ), .B(\U3/U199/Z_0 ), .Z(n5851) );
  XOR2_X1 U3788 ( .A(\U3/U196/Z_0 ), .B(\U3/U195/Z_0 ), .Z(n5852) );
  AND2_X1 U3789 ( .A1(\U3/U200/Z_0 ), .A2(\U3/U199/Z_0 ), .ZN(n5853) );
  AND2_X1 U3790 ( .A1(\U3/U200/Z_0 ), .A2(\U3/U199/Z_0 ), .ZN(n5854) );
  XOR2_X1 U3791 ( .A(\U3/U202/Z_0 ), .B(\U3/U201/Z_0 ), .Z(n5855) );
  XOR2_X1 U3792 ( .A(\U3/U200/Z_4 ), .B(\r642/carry[4] ), .Z(n5856) );
  INV_X1 U3793 ( .A(n5861), .ZN(n5865) );
  XNOR2_X1 U3794 ( .A(CWP[3]), .B(n5861), .ZN(N915) );
  XNOR2_X1 U3795 ( .A(CWP[4]), .B(\sub_128_C208/carry[4] ), .ZN(N916) );
  NAND2_X1 U3796 ( .A1(n1315), .A2(n5865), .ZN(\sub_128_C208/carry[4] ) );
  XOR2_X1 U3797 ( .A(N888), .B(ADD_WR[0]), .Z(n5857) );
  XOR2_X1 U3798 ( .A(CWP[4]), .B(\r467/carry[4] ), .Z(n5858) );
  XNOR2_X1 U3799 ( .A(CWP[2]), .B(CWP[1]), .ZN(N890) );
  XNOR2_X1 U3800 ( .A(CWP[2]), .B(CWP[1]), .ZN(n5866) );
  OR2_X1 U3801 ( .A1(CWP[2]), .A2(CWP[1]), .ZN(\r473/carry[3] ) );
  AND2_X1 U3802 ( .A1(N888), .A2(ADD_WR[0]), .ZN(n5859) );
  XOR2_X1 U3803 ( .A(\U3/U201/Z_4 ), .B(\r507/carry[4] ), .Z(n5860) );
  AND2_X1 U3804 ( .A1(CWP[2]), .A2(CWP[1]), .ZN(n5861) );
  XOR2_X1 U3805 ( .A(CWP[3]), .B(\r473/carry[3] ), .Z(n5862) );
  XOR2_X1 U3806 ( .A(n1303), .B(n5869), .Z(n5863) );
  NAND2_X1 U3807 ( .A1(CWP[3]), .A2(\r473/carry[3] ), .ZN(n5869) );
  XOR2_X1 U3808 ( .A(\U3/U196/Z_4 ), .B(\r638/carry[4] ), .Z(n5864) );
  OAI22_X1 U3809 ( .A1(n7861), .A2(n5870), .B1(n5871), .B2(n5872), .ZN(n8311)
         );
  NOR4_X1 U3810 ( .A1(n5873), .A2(n5874), .A3(n5875), .A4(n5876), .ZN(n5871)
         );
  OAI221_X1 U3811 ( .B1(n5830), .B2(n4894), .C1(n5877), .C2(n5089), .A(n5878), 
        .ZN(n5876) );
  AOI22_X1 U3812 ( .A1(n5879), .A2(n5299), .B1(n5880), .B2(n5024), .ZN(n5878)
         );
  OAI221_X1 U3813 ( .B1(n482), .B2(n5881), .C1(n546), .C2(n5882), .A(n5883), 
        .ZN(n5875) );
  AOI22_X1 U3814 ( .A1(n8053), .A2(n5884), .B1(n7989), .B2(n5885), .ZN(n5883)
         );
  OAI221_X1 U3815 ( .B1(n738), .B2(n5819), .C1(n802), .C2(n5886), .A(n5887), 
        .ZN(n5874) );
  AOI22_X1 U3816 ( .A1(n8181), .A2(n5888), .B1(n8117), .B2(n5889), .ZN(n5887)
         );
  OAI221_X1 U3817 ( .B1(n866), .B2(n5890), .C1(n930), .C2(n5891), .A(n5892), 
        .ZN(n5873) );
  AOI222_X1 U3818 ( .A1(n5893), .A2(n4958), .B1(n5894), .B2(n5217), .C1(n5895), 
        .C2(n5556), .ZN(n5892) );
  OAI22_X1 U3819 ( .A1(n7862), .A2(n5870), .B1(n5896), .B2(n5872), .ZN(n8312)
         );
  NOR4_X1 U3820 ( .A1(n5897), .A2(n5898), .A3(n5899), .A4(n5900), .ZN(n5896)
         );
  OAI221_X1 U3821 ( .B1(n5830), .B2(n4893), .C1(n5877), .C2(n5088), .A(n5901), 
        .ZN(n5900) );
  AOI22_X1 U3822 ( .A1(n5879), .A2(n5298), .B1(n5880), .B2(n5023), .ZN(n5901)
         );
  OAI221_X1 U3823 ( .B1(n483), .B2(n5881), .C1(n547), .C2(n5882), .A(n5902), 
        .ZN(n5899) );
  AOI22_X1 U3824 ( .A1(n8054), .A2(n5884), .B1(n7990), .B2(n5885), .ZN(n5902)
         );
  OAI221_X1 U3825 ( .B1(n739), .B2(n5819), .C1(n803), .C2(n5886), .A(n5903), 
        .ZN(n5898) );
  AOI22_X1 U3826 ( .A1(n8182), .A2(n5888), .B1(n8118), .B2(n5889), .ZN(n5903)
         );
  OAI221_X1 U3827 ( .B1(n867), .B2(n5890), .C1(n931), .C2(n5891), .A(n5904), 
        .ZN(n5897) );
  AOI222_X1 U3828 ( .A1(n5893), .A2(n4957), .B1(n5894), .B2(n5216), .C1(n5895), 
        .C2(n5555), .ZN(n5904) );
  OAI22_X1 U3829 ( .A1(n7863), .A2(n5870), .B1(n5905), .B2(n5872), .ZN(n8313)
         );
  NOR4_X1 U3830 ( .A1(n5906), .A2(n5907), .A3(n5908), .A4(n5909), .ZN(n5905)
         );
  OAI221_X1 U3831 ( .B1(n5830), .B2(n4892), .C1(n5877), .C2(n5087), .A(n5910), 
        .ZN(n5909) );
  AOI22_X1 U3832 ( .A1(n5879), .A2(n5297), .B1(n5880), .B2(n5022), .ZN(n5910)
         );
  OAI221_X1 U3833 ( .B1(n484), .B2(n5881), .C1(n548), .C2(n5882), .A(n5911), 
        .ZN(n5908) );
  AOI22_X1 U3834 ( .A1(n8055), .A2(n5884), .B1(n7991), .B2(n5885), .ZN(n5911)
         );
  OAI221_X1 U3835 ( .B1(n740), .B2(n5819), .C1(n804), .C2(n5886), .A(n5912), 
        .ZN(n5907) );
  AOI22_X1 U3836 ( .A1(n8183), .A2(n5888), .B1(n8119), .B2(n5889), .ZN(n5912)
         );
  OAI221_X1 U3837 ( .B1(n868), .B2(n5890), .C1(n932), .C2(n5891), .A(n5913), 
        .ZN(n5906) );
  AOI222_X1 U3838 ( .A1(n5893), .A2(n4956), .B1(n5894), .B2(n5215), .C1(n5895), 
        .C2(n5554), .ZN(n5913) );
  OAI22_X1 U3839 ( .A1(n7864), .A2(n5870), .B1(n5914), .B2(n5872), .ZN(n8314)
         );
  NOR4_X1 U3840 ( .A1(n5915), .A2(n5916), .A3(n5917), .A4(n5918), .ZN(n5914)
         );
  OAI221_X1 U3841 ( .B1(n5830), .B2(n4891), .C1(n5877), .C2(n5086), .A(n5919), 
        .ZN(n5918) );
  AOI22_X1 U3842 ( .A1(n5879), .A2(n5296), .B1(n5880), .B2(n5021), .ZN(n5919)
         );
  OAI221_X1 U3843 ( .B1(n485), .B2(n5881), .C1(n549), .C2(n5882), .A(n5920), 
        .ZN(n5917) );
  AOI22_X1 U3844 ( .A1(n8056), .A2(n5884), .B1(n7992), .B2(n5885), .ZN(n5920)
         );
  OAI221_X1 U3845 ( .B1(n741), .B2(n5819), .C1(n805), .C2(n5886), .A(n5921), 
        .ZN(n5916) );
  AOI22_X1 U3846 ( .A1(n8184), .A2(n5888), .B1(n8120), .B2(n5889), .ZN(n5921)
         );
  OAI221_X1 U3847 ( .B1(n869), .B2(n5890), .C1(n933), .C2(n5891), .A(n5922), 
        .ZN(n5915) );
  AOI222_X1 U3848 ( .A1(n5893), .A2(n4955), .B1(n5894), .B2(n5214), .C1(n5895), 
        .C2(n5553), .ZN(n5922) );
  OAI22_X1 U3849 ( .A1(n7865), .A2(n5870), .B1(n5923), .B2(n5872), .ZN(n8315)
         );
  NOR4_X1 U3850 ( .A1(n5924), .A2(n5925), .A3(n5926), .A4(n5927), .ZN(n5923)
         );
  OAI221_X1 U3851 ( .B1(n5830), .B2(n4890), .C1(n5877), .C2(n5085), .A(n5928), 
        .ZN(n5927) );
  AOI22_X1 U3852 ( .A1(n5879), .A2(n5295), .B1(n5880), .B2(n5020), .ZN(n5928)
         );
  OAI221_X1 U3853 ( .B1(n486), .B2(n5881), .C1(n550), .C2(n5882), .A(n5929), 
        .ZN(n5926) );
  AOI22_X1 U3854 ( .A1(n8057), .A2(n5884), .B1(n7993), .B2(n5885), .ZN(n5929)
         );
  OAI221_X1 U3855 ( .B1(n742), .B2(n5819), .C1(n806), .C2(n5886), .A(n5930), 
        .ZN(n5925) );
  AOI22_X1 U3856 ( .A1(n8185), .A2(n5888), .B1(n8121), .B2(n5889), .ZN(n5930)
         );
  OAI221_X1 U3857 ( .B1(n870), .B2(n5890), .C1(n934), .C2(n5891), .A(n5931), 
        .ZN(n5924) );
  AOI222_X1 U3858 ( .A1(n5893), .A2(n4954), .B1(n5894), .B2(n5213), .C1(n5895), 
        .C2(n5552), .ZN(n5931) );
  OAI22_X1 U3859 ( .A1(n7866), .A2(n5870), .B1(n5932), .B2(n5872), .ZN(n8316)
         );
  NOR4_X1 U3860 ( .A1(n5933), .A2(n5934), .A3(n5935), .A4(n5936), .ZN(n5932)
         );
  OAI221_X1 U3861 ( .B1(n5830), .B2(n4889), .C1(n5877), .C2(n5084), .A(n5937), 
        .ZN(n5936) );
  AOI22_X1 U3862 ( .A1(n5879), .A2(n5294), .B1(n5880), .B2(n5019), .ZN(n5937)
         );
  OAI221_X1 U3863 ( .B1(n487), .B2(n5881), .C1(n551), .C2(n5882), .A(n5938), 
        .ZN(n5935) );
  AOI22_X1 U3864 ( .A1(n8058), .A2(n5884), .B1(n7994), .B2(n5885), .ZN(n5938)
         );
  OAI221_X1 U3865 ( .B1(n743), .B2(n5819), .C1(n807), .C2(n5886), .A(n5939), 
        .ZN(n5934) );
  AOI22_X1 U3866 ( .A1(n8186), .A2(n5888), .B1(n8122), .B2(n5889), .ZN(n5939)
         );
  OAI221_X1 U3867 ( .B1(n871), .B2(n5890), .C1(n935), .C2(n5891), .A(n5940), 
        .ZN(n5933) );
  AOI222_X1 U3868 ( .A1(n5893), .A2(n4953), .B1(n5894), .B2(n5212), .C1(n5895), 
        .C2(n5551), .ZN(n5940) );
  OAI22_X1 U3869 ( .A1(n7867), .A2(n5870), .B1(n5941), .B2(n5872), .ZN(n8317)
         );
  NOR4_X1 U3870 ( .A1(n5942), .A2(n5943), .A3(n5944), .A4(n5945), .ZN(n5941)
         );
  OAI221_X1 U3871 ( .B1(n5830), .B2(n4888), .C1(n5877), .C2(n5083), .A(n5946), 
        .ZN(n5945) );
  AOI22_X1 U3872 ( .A1(n5879), .A2(n5293), .B1(n5880), .B2(n5018), .ZN(n5946)
         );
  OAI221_X1 U3873 ( .B1(n488), .B2(n5881), .C1(n552), .C2(n5882), .A(n5947), 
        .ZN(n5944) );
  AOI22_X1 U3874 ( .A1(n8059), .A2(n5884), .B1(n7995), .B2(n5885), .ZN(n5947)
         );
  OAI221_X1 U3875 ( .B1(n744), .B2(n5819), .C1(n808), .C2(n5886), .A(n5948), 
        .ZN(n5943) );
  AOI22_X1 U3876 ( .A1(n8187), .A2(n5888), .B1(n8123), .B2(n5889), .ZN(n5948)
         );
  OAI221_X1 U3877 ( .B1(n872), .B2(n5890), .C1(n936), .C2(n5891), .A(n5949), 
        .ZN(n5942) );
  AOI222_X1 U3878 ( .A1(n5893), .A2(n4952), .B1(n5894), .B2(n5211), .C1(n5895), 
        .C2(n5550), .ZN(n5949) );
  OAI22_X1 U3879 ( .A1(n7868), .A2(n5870), .B1(n5950), .B2(n5872), .ZN(n8318)
         );
  NOR4_X1 U3880 ( .A1(n5951), .A2(n5952), .A3(n5953), .A4(n5954), .ZN(n5950)
         );
  OAI221_X1 U3881 ( .B1(n5830), .B2(n4887), .C1(n5877), .C2(n5082), .A(n5955), 
        .ZN(n5954) );
  AOI22_X1 U3882 ( .A1(n5879), .A2(n5292), .B1(n5880), .B2(n5017), .ZN(n5955)
         );
  OAI221_X1 U3883 ( .B1(n489), .B2(n5881), .C1(n553), .C2(n5882), .A(n5956), 
        .ZN(n5953) );
  AOI22_X1 U3884 ( .A1(n8060), .A2(n5884), .B1(n7996), .B2(n5885), .ZN(n5956)
         );
  OAI221_X1 U3885 ( .B1(n745), .B2(n5819), .C1(n809), .C2(n5886), .A(n5957), 
        .ZN(n5952) );
  AOI22_X1 U3886 ( .A1(n8188), .A2(n5888), .B1(n8124), .B2(n5889), .ZN(n5957)
         );
  OAI221_X1 U3887 ( .B1(n873), .B2(n5890), .C1(n937), .C2(n5891), .A(n5958), 
        .ZN(n5951) );
  AOI222_X1 U3888 ( .A1(n5893), .A2(n4951), .B1(n5894), .B2(n5210), .C1(n5895), 
        .C2(n5549), .ZN(n5958) );
  OAI22_X1 U3889 ( .A1(n7869), .A2(n5870), .B1(n5959), .B2(n5872), .ZN(n8319)
         );
  NOR4_X1 U3890 ( .A1(n5960), .A2(n5961), .A3(n5962), .A4(n5963), .ZN(n5959)
         );
  OAI221_X1 U3891 ( .B1(n5830), .B2(n4886), .C1(n5877), .C2(n5081), .A(n5964), 
        .ZN(n5963) );
  AOI22_X1 U3892 ( .A1(n5879), .A2(n5291), .B1(n5880), .B2(n5016), .ZN(n5964)
         );
  OAI221_X1 U3893 ( .B1(n490), .B2(n5881), .C1(n554), .C2(n5882), .A(n5965), 
        .ZN(n5962) );
  AOI22_X1 U3894 ( .A1(n8061), .A2(n5884), .B1(n7997), .B2(n5885), .ZN(n5965)
         );
  OAI221_X1 U3895 ( .B1(n746), .B2(n5819), .C1(n810), .C2(n5886), .A(n5966), 
        .ZN(n5961) );
  AOI22_X1 U3896 ( .A1(n8189), .A2(n5888), .B1(n8125), .B2(n5889), .ZN(n5966)
         );
  OAI221_X1 U3897 ( .B1(n874), .B2(n5890), .C1(n938), .C2(n5891), .A(n5967), 
        .ZN(n5960) );
  AOI222_X1 U3898 ( .A1(n5893), .A2(n4950), .B1(n5894), .B2(n5209), .C1(n5895), 
        .C2(n5548), .ZN(n5967) );
  OAI22_X1 U3899 ( .A1(n7870), .A2(n5870), .B1(n5968), .B2(n5872), .ZN(n8320)
         );
  NOR4_X1 U3900 ( .A1(n5969), .A2(n5970), .A3(n5971), .A4(n5972), .ZN(n5968)
         );
  OAI221_X1 U3901 ( .B1(n5830), .B2(n4885), .C1(n5877), .C2(n5080), .A(n5973), 
        .ZN(n5972) );
  AOI22_X1 U3902 ( .A1(n5879), .A2(n5290), .B1(n5880), .B2(n5015), .ZN(n5973)
         );
  OAI221_X1 U3903 ( .B1(n491), .B2(n5881), .C1(n555), .C2(n5882), .A(n5974), 
        .ZN(n5971) );
  AOI22_X1 U3904 ( .A1(n8062), .A2(n5884), .B1(n7998), .B2(n5885), .ZN(n5974)
         );
  OAI221_X1 U3905 ( .B1(n747), .B2(n5819), .C1(n811), .C2(n5886), .A(n5975), 
        .ZN(n5970) );
  AOI22_X1 U3906 ( .A1(n8190), .A2(n5888), .B1(n8126), .B2(n5889), .ZN(n5975)
         );
  OAI221_X1 U3907 ( .B1(n875), .B2(n5890), .C1(n939), .C2(n5891), .A(n5976), 
        .ZN(n5969) );
  AOI222_X1 U3908 ( .A1(n5893), .A2(n4949), .B1(n5894), .B2(n5208), .C1(n5895), 
        .C2(n5547), .ZN(n5976) );
  OAI22_X1 U3909 ( .A1(n7871), .A2(n5870), .B1(n5977), .B2(n5872), .ZN(n8321)
         );
  NOR4_X1 U3910 ( .A1(n5978), .A2(n5979), .A3(n5980), .A4(n5981), .ZN(n5977)
         );
  OAI221_X1 U3911 ( .B1(n5830), .B2(n4884), .C1(n5877), .C2(n5079), .A(n5982), 
        .ZN(n5981) );
  AOI22_X1 U3912 ( .A1(n5879), .A2(n5289), .B1(n5880), .B2(n5014), .ZN(n5982)
         );
  OAI221_X1 U3913 ( .B1(n492), .B2(n5881), .C1(n556), .C2(n5882), .A(n5983), 
        .ZN(n5980) );
  AOI22_X1 U3914 ( .A1(n8063), .A2(n5884), .B1(n7999), .B2(n5885), .ZN(n5983)
         );
  OAI221_X1 U3915 ( .B1(n748), .B2(n5819), .C1(n812), .C2(n5886), .A(n5984), 
        .ZN(n5979) );
  AOI22_X1 U3916 ( .A1(n8191), .A2(n5888), .B1(n8127), .B2(n5889), .ZN(n5984)
         );
  OAI221_X1 U3917 ( .B1(n876), .B2(n5890), .C1(n940), .C2(n5891), .A(n5985), 
        .ZN(n5978) );
  AOI222_X1 U3918 ( .A1(n5893), .A2(n4948), .B1(n5894), .B2(n5207), .C1(n5895), 
        .C2(n5546), .ZN(n5985) );
  OAI22_X1 U3919 ( .A1(n7872), .A2(n5870), .B1(n5986), .B2(n5872), .ZN(n8322)
         );
  NOR4_X1 U3920 ( .A1(n5987), .A2(n5988), .A3(n5989), .A4(n5990), .ZN(n5986)
         );
  OAI221_X1 U3921 ( .B1(n5830), .B2(n4883), .C1(n5877), .C2(n5078), .A(n5991), 
        .ZN(n5990) );
  AOI22_X1 U3922 ( .A1(n5879), .A2(n5288), .B1(n5880), .B2(n5013), .ZN(n5991)
         );
  OAI221_X1 U3923 ( .B1(n493), .B2(n5881), .C1(n557), .C2(n5882), .A(n5992), 
        .ZN(n5989) );
  AOI22_X1 U3924 ( .A1(n8064), .A2(n5884), .B1(n8000), .B2(n5885), .ZN(n5992)
         );
  OAI221_X1 U3925 ( .B1(n749), .B2(n5819), .C1(n813), .C2(n5886), .A(n5993), 
        .ZN(n5988) );
  AOI22_X1 U3926 ( .A1(n8192), .A2(n5888), .B1(n8128), .B2(n5889), .ZN(n5993)
         );
  OAI221_X1 U3927 ( .B1(n877), .B2(n5890), .C1(n941), .C2(n5891), .A(n5994), 
        .ZN(n5987) );
  AOI222_X1 U3928 ( .A1(n5893), .A2(n4947), .B1(n5894), .B2(n5206), .C1(n5895), 
        .C2(n5545), .ZN(n5994) );
  OAI22_X1 U3929 ( .A1(n7873), .A2(n5870), .B1(n5995), .B2(n5872), .ZN(n8323)
         );
  NOR4_X1 U3930 ( .A1(n5996), .A2(n5997), .A3(n5998), .A4(n5999), .ZN(n5995)
         );
  OAI221_X1 U3931 ( .B1(n5830), .B2(n4882), .C1(n5877), .C2(n5077), .A(n6000), 
        .ZN(n5999) );
  AOI22_X1 U3932 ( .A1(n5879), .A2(n5287), .B1(n5880), .B2(n5012), .ZN(n6000)
         );
  OAI221_X1 U3933 ( .B1(n494), .B2(n5881), .C1(n558), .C2(n5882), .A(n6001), 
        .ZN(n5998) );
  AOI22_X1 U3934 ( .A1(n8065), .A2(n5884), .B1(n8001), .B2(n5885), .ZN(n6001)
         );
  OAI221_X1 U3935 ( .B1(n750), .B2(n5819), .C1(n814), .C2(n5886), .A(n6002), 
        .ZN(n5997) );
  AOI22_X1 U3936 ( .A1(n8193), .A2(n5888), .B1(n8129), .B2(n5889), .ZN(n6002)
         );
  OAI221_X1 U3937 ( .B1(n878), .B2(n5890), .C1(n942), .C2(n5891), .A(n6003), 
        .ZN(n5996) );
  AOI222_X1 U3938 ( .A1(n5893), .A2(n4946), .B1(n5894), .B2(n5205), .C1(n5895), 
        .C2(n5544), .ZN(n6003) );
  OAI22_X1 U3939 ( .A1(n7874), .A2(n5870), .B1(n6004), .B2(n5872), .ZN(n8324)
         );
  NOR4_X1 U3940 ( .A1(n6005), .A2(n6006), .A3(n6007), .A4(n6008), .ZN(n6004)
         );
  OAI221_X1 U3941 ( .B1(n5830), .B2(n4881), .C1(n5877), .C2(n5076), .A(n6009), 
        .ZN(n6008) );
  AOI22_X1 U3942 ( .A1(n5879), .A2(n5286), .B1(n5880), .B2(n5011), .ZN(n6009)
         );
  OAI221_X1 U3943 ( .B1(n495), .B2(n5881), .C1(n559), .C2(n5882), .A(n6010), 
        .ZN(n6007) );
  AOI22_X1 U3944 ( .A1(n8066), .A2(n5884), .B1(n8002), .B2(n5885), .ZN(n6010)
         );
  OAI221_X1 U3945 ( .B1(n751), .B2(n5819), .C1(n815), .C2(n5886), .A(n6011), 
        .ZN(n6006) );
  AOI22_X1 U3946 ( .A1(n8194), .A2(n5888), .B1(n8130), .B2(n5889), .ZN(n6011)
         );
  OAI221_X1 U3947 ( .B1(n879), .B2(n5890), .C1(n943), .C2(n5891), .A(n6012), 
        .ZN(n6005) );
  AOI222_X1 U3948 ( .A1(n5893), .A2(n4945), .B1(n5894), .B2(n5204), .C1(n5895), 
        .C2(n5543), .ZN(n6012) );
  OAI22_X1 U3949 ( .A1(n7875), .A2(n5870), .B1(n6013), .B2(n5872), .ZN(n8325)
         );
  NOR4_X1 U3950 ( .A1(n6014), .A2(n6015), .A3(n6016), .A4(n6017), .ZN(n6013)
         );
  OAI221_X1 U3951 ( .B1(n5830), .B2(n4880), .C1(n5877), .C2(n5075), .A(n6018), 
        .ZN(n6017) );
  AOI22_X1 U3952 ( .A1(n5879), .A2(n5285), .B1(n5880), .B2(n5010), .ZN(n6018)
         );
  OAI221_X1 U3953 ( .B1(n496), .B2(n5881), .C1(n560), .C2(n5882), .A(n6019), 
        .ZN(n6016) );
  AOI22_X1 U3954 ( .A1(n8067), .A2(n5884), .B1(n8003), .B2(n5885), .ZN(n6019)
         );
  OAI221_X1 U3955 ( .B1(n752), .B2(n5819), .C1(n816), .C2(n5886), .A(n6020), 
        .ZN(n6015) );
  AOI22_X1 U3956 ( .A1(n8195), .A2(n5888), .B1(n8131), .B2(n5889), .ZN(n6020)
         );
  OAI221_X1 U3957 ( .B1(n880), .B2(n5890), .C1(n944), .C2(n5891), .A(n6021), 
        .ZN(n6014) );
  AOI222_X1 U3958 ( .A1(n5893), .A2(n4944), .B1(n5894), .B2(n5203), .C1(n5895), 
        .C2(n5542), .ZN(n6021) );
  OAI22_X1 U3959 ( .A1(n7876), .A2(n5870), .B1(n6022), .B2(n5872), .ZN(n8326)
         );
  NOR4_X1 U3960 ( .A1(n6023), .A2(n6024), .A3(n6025), .A4(n6026), .ZN(n6022)
         );
  OAI221_X1 U3961 ( .B1(n5830), .B2(n4879), .C1(n5877), .C2(n5074), .A(n6027), 
        .ZN(n6026) );
  AOI22_X1 U3962 ( .A1(n5879), .A2(n5284), .B1(n5880), .B2(n5009), .ZN(n6027)
         );
  OAI221_X1 U3963 ( .B1(n497), .B2(n5881), .C1(n561), .C2(n5882), .A(n6028), 
        .ZN(n6025) );
  AOI22_X1 U3964 ( .A1(n8068), .A2(n5884), .B1(n8004), .B2(n5885), .ZN(n6028)
         );
  OAI221_X1 U3965 ( .B1(n753), .B2(n5819), .C1(n817), .C2(n5886), .A(n6029), 
        .ZN(n6024) );
  AOI22_X1 U3966 ( .A1(n8196), .A2(n5888), .B1(n8132), .B2(n5889), .ZN(n6029)
         );
  OAI221_X1 U3967 ( .B1(n881), .B2(n5890), .C1(n945), .C2(n5891), .A(n6030), 
        .ZN(n6023) );
  AOI222_X1 U3968 ( .A1(n5893), .A2(n4943), .B1(n5894), .B2(n5202), .C1(n5895), 
        .C2(n5541), .ZN(n6030) );
  OAI22_X1 U3969 ( .A1(n7877), .A2(n5870), .B1(n6031), .B2(n5872), .ZN(n8327)
         );
  NOR4_X1 U3970 ( .A1(n6032), .A2(n6033), .A3(n6034), .A4(n6035), .ZN(n6031)
         );
  OAI221_X1 U3971 ( .B1(n5830), .B2(n4878), .C1(n5877), .C2(n5073), .A(n6036), 
        .ZN(n6035) );
  AOI22_X1 U3972 ( .A1(n5879), .A2(n5283), .B1(n5880), .B2(n5008), .ZN(n6036)
         );
  OAI221_X1 U3973 ( .B1(n498), .B2(n5881), .C1(n562), .C2(n5882), .A(n6037), 
        .ZN(n6034) );
  AOI22_X1 U3974 ( .A1(n8069), .A2(n5884), .B1(n8005), .B2(n5885), .ZN(n6037)
         );
  OAI221_X1 U3975 ( .B1(n754), .B2(n5819), .C1(n818), .C2(n5886), .A(n6038), 
        .ZN(n6033) );
  AOI22_X1 U3976 ( .A1(n8197), .A2(n5888), .B1(n8133), .B2(n5889), .ZN(n6038)
         );
  OAI221_X1 U3977 ( .B1(n882), .B2(n5890), .C1(n946), .C2(n5891), .A(n6039), 
        .ZN(n6032) );
  AOI222_X1 U3978 ( .A1(n5893), .A2(n4942), .B1(n5894), .B2(n5201), .C1(n5895), 
        .C2(n5540), .ZN(n6039) );
  OAI22_X1 U3979 ( .A1(n7878), .A2(n5870), .B1(n6040), .B2(n5872), .ZN(n8328)
         );
  NOR4_X1 U3980 ( .A1(n6041), .A2(n6042), .A3(n6043), .A4(n6044), .ZN(n6040)
         );
  OAI221_X1 U3981 ( .B1(n5830), .B2(n4877), .C1(n5877), .C2(n5072), .A(n6045), 
        .ZN(n6044) );
  AOI22_X1 U3982 ( .A1(n5879), .A2(n5282), .B1(n5880), .B2(n5007), .ZN(n6045)
         );
  OAI221_X1 U3983 ( .B1(n499), .B2(n5881), .C1(n563), .C2(n5882), .A(n6046), 
        .ZN(n6043) );
  AOI22_X1 U3984 ( .A1(n8070), .A2(n5884), .B1(n8006), .B2(n5885), .ZN(n6046)
         );
  OAI221_X1 U3985 ( .B1(n755), .B2(n5819), .C1(n819), .C2(n5886), .A(n6047), 
        .ZN(n6042) );
  AOI22_X1 U3986 ( .A1(n8198), .A2(n5888), .B1(n8134), .B2(n5889), .ZN(n6047)
         );
  OAI221_X1 U3987 ( .B1(n883), .B2(n5890), .C1(n947), .C2(n5891), .A(n6048), 
        .ZN(n6041) );
  AOI222_X1 U3988 ( .A1(n5893), .A2(n4941), .B1(n5894), .B2(n5200), .C1(n5895), 
        .C2(n5539), .ZN(n6048) );
  OAI22_X1 U3989 ( .A1(n7879), .A2(n5870), .B1(n6049), .B2(n5872), .ZN(n8329)
         );
  NOR4_X1 U3990 ( .A1(n6050), .A2(n6051), .A3(n6052), .A4(n6053), .ZN(n6049)
         );
  OAI221_X1 U3991 ( .B1(n5830), .B2(n4876), .C1(n5877), .C2(n5071), .A(n6054), 
        .ZN(n6053) );
  AOI22_X1 U3992 ( .A1(n5879), .A2(n5281), .B1(n5880), .B2(n5006), .ZN(n6054)
         );
  OAI221_X1 U3993 ( .B1(n500), .B2(n5881), .C1(n564), .C2(n5882), .A(n6055), 
        .ZN(n6052) );
  AOI22_X1 U3994 ( .A1(n8071), .A2(n5884), .B1(n8007), .B2(n5885), .ZN(n6055)
         );
  OAI221_X1 U3995 ( .B1(n756), .B2(n5819), .C1(n820), .C2(n5886), .A(n6056), 
        .ZN(n6051) );
  AOI22_X1 U3996 ( .A1(n8199), .A2(n5888), .B1(n8135), .B2(n5889), .ZN(n6056)
         );
  OAI221_X1 U3997 ( .B1(n884), .B2(n5890), .C1(n948), .C2(n5891), .A(n6057), 
        .ZN(n6050) );
  AOI222_X1 U3998 ( .A1(n5893), .A2(n4940), .B1(n5894), .B2(n5199), .C1(n5895), 
        .C2(n5538), .ZN(n6057) );
  OAI22_X1 U3999 ( .A1(n7880), .A2(n5870), .B1(n6058), .B2(n5872), .ZN(n8330)
         );
  NOR4_X1 U4000 ( .A1(n6059), .A2(n6060), .A3(n6061), .A4(n6062), .ZN(n6058)
         );
  OAI221_X1 U4001 ( .B1(n5830), .B2(n4875), .C1(n5877), .C2(n5070), .A(n6063), 
        .ZN(n6062) );
  AOI22_X1 U4002 ( .A1(n5879), .A2(n5280), .B1(n5880), .B2(n5005), .ZN(n6063)
         );
  OAI221_X1 U4003 ( .B1(n501), .B2(n5881), .C1(n565), .C2(n5882), .A(n6064), 
        .ZN(n6061) );
  AOI22_X1 U4004 ( .A1(n8072), .A2(n5884), .B1(n8008), .B2(n5885), .ZN(n6064)
         );
  OAI221_X1 U4005 ( .B1(n757), .B2(n5819), .C1(n821), .C2(n5886), .A(n6065), 
        .ZN(n6060) );
  AOI22_X1 U4006 ( .A1(n8200), .A2(n5888), .B1(n8136), .B2(n5889), .ZN(n6065)
         );
  OAI221_X1 U4007 ( .B1(n885), .B2(n5890), .C1(n949), .C2(n5891), .A(n6066), 
        .ZN(n6059) );
  AOI222_X1 U4008 ( .A1(n5893), .A2(n4939), .B1(n5894), .B2(n5198), .C1(n5895), 
        .C2(n5537), .ZN(n6066) );
  OAI22_X1 U4009 ( .A1(n7881), .A2(n5870), .B1(n6067), .B2(n5872), .ZN(n8331)
         );
  NOR4_X1 U4010 ( .A1(n6068), .A2(n6069), .A3(n6070), .A4(n6071), .ZN(n6067)
         );
  OAI221_X1 U4011 ( .B1(n5830), .B2(n4874), .C1(n5877), .C2(n5069), .A(n6072), 
        .ZN(n6071) );
  AOI22_X1 U4012 ( .A1(n5879), .A2(n5279), .B1(n5880), .B2(n5004), .ZN(n6072)
         );
  OAI221_X1 U4013 ( .B1(n502), .B2(n5881), .C1(n566), .C2(n5882), .A(n6073), 
        .ZN(n6070) );
  AOI22_X1 U4014 ( .A1(n8073), .A2(n5884), .B1(n8009), .B2(n5885), .ZN(n6073)
         );
  OAI221_X1 U4015 ( .B1(n758), .B2(n5819), .C1(n822), .C2(n5886), .A(n6074), 
        .ZN(n6069) );
  AOI22_X1 U4016 ( .A1(n8201), .A2(n5888), .B1(n8137), .B2(n5889), .ZN(n6074)
         );
  OAI221_X1 U4017 ( .B1(n886), .B2(n5890), .C1(n950), .C2(n5891), .A(n6075), 
        .ZN(n6068) );
  AOI222_X1 U4018 ( .A1(n5893), .A2(n4938), .B1(n5894), .B2(n5197), .C1(n5895), 
        .C2(n5536), .ZN(n6075) );
  OAI22_X1 U4019 ( .A1(n7882), .A2(n5870), .B1(n6076), .B2(n5872), .ZN(n8332)
         );
  NOR4_X1 U4020 ( .A1(n6077), .A2(n6078), .A3(n6079), .A4(n6080), .ZN(n6076)
         );
  OAI221_X1 U4021 ( .B1(n5830), .B2(n4873), .C1(n5877), .C2(n5068), .A(n6081), 
        .ZN(n6080) );
  AOI22_X1 U4022 ( .A1(n5879), .A2(n5278), .B1(n5880), .B2(n5003), .ZN(n6081)
         );
  OAI221_X1 U4023 ( .B1(n503), .B2(n5881), .C1(n567), .C2(n5882), .A(n6082), 
        .ZN(n6079) );
  AOI22_X1 U4024 ( .A1(n8074), .A2(n5884), .B1(n8010), .B2(n5885), .ZN(n6082)
         );
  OAI221_X1 U4025 ( .B1(n759), .B2(n5819), .C1(n823), .C2(n5886), .A(n6083), 
        .ZN(n6078) );
  AOI22_X1 U4026 ( .A1(n8202), .A2(n5888), .B1(n8138), .B2(n5889), .ZN(n6083)
         );
  OAI221_X1 U4027 ( .B1(n887), .B2(n5890), .C1(n951), .C2(n5891), .A(n6084), 
        .ZN(n6077) );
  AOI222_X1 U4028 ( .A1(n5893), .A2(n4937), .B1(n5894), .B2(n5196), .C1(n5895), 
        .C2(n5535), .ZN(n6084) );
  OAI22_X1 U4029 ( .A1(n7883), .A2(n5870), .B1(n6085), .B2(n5872), .ZN(n8333)
         );
  NOR4_X1 U4030 ( .A1(n6086), .A2(n6087), .A3(n6088), .A4(n6089), .ZN(n6085)
         );
  OAI221_X1 U4031 ( .B1(n5830), .B2(n4872), .C1(n5877), .C2(n5067), .A(n6090), 
        .ZN(n6089) );
  AOI22_X1 U4032 ( .A1(n5879), .A2(n5277), .B1(n5880), .B2(n5002), .ZN(n6090)
         );
  OAI221_X1 U4033 ( .B1(n504), .B2(n5881), .C1(n568), .C2(n5882), .A(n6091), 
        .ZN(n6088) );
  AOI22_X1 U4034 ( .A1(n8075), .A2(n5884), .B1(n8011), .B2(n5885), .ZN(n6091)
         );
  OAI221_X1 U4035 ( .B1(n760), .B2(n5819), .C1(n824), .C2(n5886), .A(n6092), 
        .ZN(n6087) );
  AOI22_X1 U4036 ( .A1(n8203), .A2(n5888), .B1(n8139), .B2(n5889), .ZN(n6092)
         );
  OAI221_X1 U4037 ( .B1(n888), .B2(n5890), .C1(n952), .C2(n5891), .A(n6093), 
        .ZN(n6086) );
  AOI222_X1 U4038 ( .A1(n5893), .A2(n4936), .B1(n5894), .B2(n5195), .C1(n5895), 
        .C2(n5534), .ZN(n6093) );
  OAI22_X1 U4039 ( .A1(n7884), .A2(n5870), .B1(n6094), .B2(n5872), .ZN(n8334)
         );
  NOR4_X1 U4040 ( .A1(n6095), .A2(n6096), .A3(n6097), .A4(n6098), .ZN(n6094)
         );
  OAI221_X1 U4041 ( .B1(n5830), .B2(n4871), .C1(n5877), .C2(n5066), .A(n6099), 
        .ZN(n6098) );
  AOI22_X1 U4042 ( .A1(n5879), .A2(n5276), .B1(n5880), .B2(n5001), .ZN(n6099)
         );
  OAI221_X1 U4043 ( .B1(n505), .B2(n5881), .C1(n569), .C2(n5882), .A(n6100), 
        .ZN(n6097) );
  AOI22_X1 U4044 ( .A1(n8076), .A2(n5884), .B1(n8012), .B2(n5885), .ZN(n6100)
         );
  OAI221_X1 U4045 ( .B1(n761), .B2(n5819), .C1(n825), .C2(n5886), .A(n6101), 
        .ZN(n6096) );
  AOI22_X1 U4046 ( .A1(n8204), .A2(n5888), .B1(n8140), .B2(n5889), .ZN(n6101)
         );
  OAI221_X1 U4047 ( .B1(n889), .B2(n5890), .C1(n953), .C2(n5891), .A(n6102), 
        .ZN(n6095) );
  AOI222_X1 U4048 ( .A1(n5893), .A2(n4935), .B1(n5894), .B2(n5194), .C1(n5895), 
        .C2(n5533), .ZN(n6102) );
  OAI22_X1 U4049 ( .A1(n7885), .A2(n5870), .B1(n6103), .B2(n5872), .ZN(n8335)
         );
  NOR4_X1 U4050 ( .A1(n6104), .A2(n6105), .A3(n6106), .A4(n6107), .ZN(n6103)
         );
  OAI221_X1 U4051 ( .B1(n5830), .B2(n4870), .C1(n5877), .C2(n5065), .A(n6108), 
        .ZN(n6107) );
  AOI22_X1 U4052 ( .A1(n5879), .A2(n5275), .B1(n5880), .B2(n5000), .ZN(n6108)
         );
  OAI221_X1 U4053 ( .B1(n506), .B2(n5881), .C1(n570), .C2(n5882), .A(n6109), 
        .ZN(n6106) );
  AOI22_X1 U4054 ( .A1(n8077), .A2(n5884), .B1(n8013), .B2(n5885), .ZN(n6109)
         );
  OAI221_X1 U4055 ( .B1(n762), .B2(n5819), .C1(n826), .C2(n5886), .A(n6110), 
        .ZN(n6105) );
  AOI22_X1 U4056 ( .A1(n8205), .A2(n5888), .B1(n8141), .B2(n5889), .ZN(n6110)
         );
  OAI221_X1 U4057 ( .B1(n890), .B2(n5890), .C1(n954), .C2(n5891), .A(n6111), 
        .ZN(n6104) );
  AOI222_X1 U4058 ( .A1(n5893), .A2(n4934), .B1(n5894), .B2(n5193), .C1(n5895), 
        .C2(n5532), .ZN(n6111) );
  OAI22_X1 U4059 ( .A1(n7886), .A2(n5870), .B1(n6112), .B2(n5872), .ZN(n8336)
         );
  NOR4_X1 U4060 ( .A1(n6113), .A2(n6114), .A3(n6115), .A4(n6116), .ZN(n6112)
         );
  OAI221_X1 U4061 ( .B1(n5830), .B2(n4869), .C1(n5877), .C2(n5064), .A(n6117), 
        .ZN(n6116) );
  AOI22_X1 U4062 ( .A1(n5879), .A2(n5274), .B1(n5880), .B2(n4999), .ZN(n6117)
         );
  OAI221_X1 U4063 ( .B1(n507), .B2(n5881), .C1(n571), .C2(n5882), .A(n6118), 
        .ZN(n6115) );
  AOI22_X1 U4064 ( .A1(n8078), .A2(n5884), .B1(n8014), .B2(n5885), .ZN(n6118)
         );
  OAI221_X1 U4065 ( .B1(n763), .B2(n5819), .C1(n827), .C2(n5886), .A(n6119), 
        .ZN(n6114) );
  AOI22_X1 U4066 ( .A1(n8206), .A2(n5888), .B1(n8142), .B2(n5889), .ZN(n6119)
         );
  OAI221_X1 U4067 ( .B1(n891), .B2(n5890), .C1(n955), .C2(n5891), .A(n6120), 
        .ZN(n6113) );
  AOI222_X1 U4068 ( .A1(n5893), .A2(n4933), .B1(n5894), .B2(n5192), .C1(n5895), 
        .C2(n5531), .ZN(n6120) );
  OAI22_X1 U4069 ( .A1(n7887), .A2(n5870), .B1(n6121), .B2(n5872), .ZN(n8337)
         );
  NOR4_X1 U4070 ( .A1(n6122), .A2(n6123), .A3(n6124), .A4(n6125), .ZN(n6121)
         );
  OAI221_X1 U4071 ( .B1(n5830), .B2(n4868), .C1(n5877), .C2(n5063), .A(n6126), 
        .ZN(n6125) );
  AOI22_X1 U4072 ( .A1(n5879), .A2(n5273), .B1(n5880), .B2(n4998), .ZN(n6126)
         );
  OAI221_X1 U4073 ( .B1(n508), .B2(n5881), .C1(n572), .C2(n5882), .A(n6127), 
        .ZN(n6124) );
  AOI22_X1 U4074 ( .A1(n8079), .A2(n5884), .B1(n8015), .B2(n5885), .ZN(n6127)
         );
  OAI221_X1 U4075 ( .B1(n764), .B2(n5819), .C1(n828), .C2(n5886), .A(n6128), 
        .ZN(n6123) );
  AOI22_X1 U4076 ( .A1(n8207), .A2(n5888), .B1(n8143), .B2(n5889), .ZN(n6128)
         );
  OAI221_X1 U4077 ( .B1(n892), .B2(n5890), .C1(n956), .C2(n5891), .A(n6129), 
        .ZN(n6122) );
  AOI222_X1 U4078 ( .A1(n5893), .A2(n4932), .B1(n5894), .B2(n5191), .C1(n5895), 
        .C2(n5530), .ZN(n6129) );
  OAI22_X1 U4079 ( .A1(n7888), .A2(n5870), .B1(n6130), .B2(n5872), .ZN(n8338)
         );
  NOR4_X1 U4080 ( .A1(n6131), .A2(n6132), .A3(n6133), .A4(n6134), .ZN(n6130)
         );
  OAI221_X1 U4081 ( .B1(n5830), .B2(n4867), .C1(n5877), .C2(n5062), .A(n6135), 
        .ZN(n6134) );
  AOI22_X1 U4082 ( .A1(n5879), .A2(n5272), .B1(n5880), .B2(n4997), .ZN(n6135)
         );
  OAI221_X1 U4083 ( .B1(n509), .B2(n5881), .C1(n573), .C2(n5882), .A(n6136), 
        .ZN(n6133) );
  AOI22_X1 U4084 ( .A1(n8080), .A2(n5884), .B1(n8016), .B2(n5885), .ZN(n6136)
         );
  OAI221_X1 U4085 ( .B1(n765), .B2(n5819), .C1(n829), .C2(n5886), .A(n6137), 
        .ZN(n6132) );
  AOI22_X1 U4086 ( .A1(n8208), .A2(n5888), .B1(n8144), .B2(n5889), .ZN(n6137)
         );
  OAI221_X1 U4087 ( .B1(n893), .B2(n5890), .C1(n957), .C2(n5891), .A(n6138), 
        .ZN(n6131) );
  AOI222_X1 U4088 ( .A1(n5893), .A2(n4931), .B1(n5894), .B2(n5190), .C1(n5895), 
        .C2(n5529), .ZN(n6138) );
  OAI22_X1 U4089 ( .A1(n7889), .A2(n5870), .B1(n6139), .B2(n5872), .ZN(n8339)
         );
  NOR4_X1 U4090 ( .A1(n6140), .A2(n6141), .A3(n6142), .A4(n6143), .ZN(n6139)
         );
  OAI221_X1 U4091 ( .B1(n5830), .B2(n4866), .C1(n5877), .C2(n5061), .A(n6144), 
        .ZN(n6143) );
  AOI22_X1 U4092 ( .A1(n5879), .A2(n5271), .B1(n5880), .B2(n4996), .ZN(n6144)
         );
  OAI221_X1 U4093 ( .B1(n510), .B2(n5881), .C1(n574), .C2(n5882), .A(n6145), 
        .ZN(n6142) );
  AOI22_X1 U4094 ( .A1(n8081), .A2(n5884), .B1(n8017), .B2(n5885), .ZN(n6145)
         );
  OAI221_X1 U4095 ( .B1(n766), .B2(n5819), .C1(n830), .C2(n5886), .A(n6146), 
        .ZN(n6141) );
  AOI22_X1 U4096 ( .A1(n8209), .A2(n5888), .B1(n8145), .B2(n5889), .ZN(n6146)
         );
  OAI221_X1 U4097 ( .B1(n894), .B2(n5890), .C1(n958), .C2(n5891), .A(n6147), 
        .ZN(n6140) );
  AOI222_X1 U4098 ( .A1(n5893), .A2(n4930), .B1(n5894), .B2(n5189), .C1(n5895), 
        .C2(n5528), .ZN(n6147) );
  OAI22_X1 U4099 ( .A1(n7890), .A2(n5870), .B1(n6148), .B2(n5872), .ZN(n8340)
         );
  NOR4_X1 U4100 ( .A1(n6149), .A2(n6150), .A3(n6151), .A4(n6152), .ZN(n6148)
         );
  OAI221_X1 U4101 ( .B1(n5830), .B2(n4865), .C1(n5877), .C2(n5060), .A(n6153), 
        .ZN(n6152) );
  AOI22_X1 U4102 ( .A1(n5879), .A2(n5270), .B1(n5880), .B2(n4995), .ZN(n6153)
         );
  OAI221_X1 U4103 ( .B1(n511), .B2(n5881), .C1(n575), .C2(n5882), .A(n6154), 
        .ZN(n6151) );
  AOI22_X1 U4104 ( .A1(n8082), .A2(n5884), .B1(n8018), .B2(n5885), .ZN(n6154)
         );
  OAI221_X1 U4105 ( .B1(n767), .B2(n5819), .C1(n831), .C2(n5886), .A(n6155), 
        .ZN(n6150) );
  AOI22_X1 U4106 ( .A1(n8210), .A2(n5888), .B1(n8146), .B2(n5889), .ZN(n6155)
         );
  OAI221_X1 U4107 ( .B1(n895), .B2(n5890), .C1(n959), .C2(n5891), .A(n6156), 
        .ZN(n6149) );
  AOI222_X1 U4108 ( .A1(n5893), .A2(n4929), .B1(n5894), .B2(n5188), .C1(n5895), 
        .C2(n5527), .ZN(n6156) );
  OAI22_X1 U4109 ( .A1(n7891), .A2(n5870), .B1(n6157), .B2(n5872), .ZN(n8341)
         );
  NOR4_X1 U4110 ( .A1(n6158), .A2(n6159), .A3(n6160), .A4(n6161), .ZN(n6157)
         );
  OAI221_X1 U4111 ( .B1(n5830), .B2(n4864), .C1(n5877), .C2(n5059), .A(n6162), 
        .ZN(n6161) );
  AOI22_X1 U4112 ( .A1(n5879), .A2(n5269), .B1(n5880), .B2(n4994), .ZN(n6162)
         );
  OAI221_X1 U4113 ( .B1(n512), .B2(n5881), .C1(n576), .C2(n5882), .A(n6163), 
        .ZN(n6160) );
  AOI22_X1 U4114 ( .A1(n8083), .A2(n5884), .B1(n8019), .B2(n5885), .ZN(n6163)
         );
  OAI221_X1 U4115 ( .B1(n768), .B2(n5819), .C1(n832), .C2(n5886), .A(n6164), 
        .ZN(n6159) );
  AOI22_X1 U4116 ( .A1(n8211), .A2(n5888), .B1(n8147), .B2(n5889), .ZN(n6164)
         );
  OAI221_X1 U4117 ( .B1(n896), .B2(n5890), .C1(n960), .C2(n5891), .A(n6165), 
        .ZN(n6158) );
  AOI222_X1 U4118 ( .A1(n5893), .A2(n4928), .B1(n5894), .B2(n5187), .C1(n5895), 
        .C2(n5526), .ZN(n6165) );
  OAI22_X1 U4119 ( .A1(n7892), .A2(n5870), .B1(n6166), .B2(n5872), .ZN(n8342)
         );
  NOR4_X1 U4120 ( .A1(n6167), .A2(n6168), .A3(n6169), .A4(n6170), .ZN(n6166)
         );
  OAI221_X1 U4121 ( .B1(n5830), .B2(n4863), .C1(n5877), .C2(n5058), .A(n6171), 
        .ZN(n6170) );
  AOI22_X1 U4122 ( .A1(n5879), .A2(n5268), .B1(n5880), .B2(n4993), .ZN(n6171)
         );
  OAI221_X1 U4123 ( .B1(n513), .B2(n5881), .C1(n577), .C2(n5882), .A(n6172), 
        .ZN(n6169) );
  AOI22_X1 U4124 ( .A1(n8084), .A2(n5884), .B1(n8020), .B2(n5885), .ZN(n6172)
         );
  OAI221_X1 U4125 ( .B1(n769), .B2(n5819), .C1(n833), .C2(n5886), .A(n6173), 
        .ZN(n6168) );
  AOI22_X1 U4126 ( .A1(n8212), .A2(n5888), .B1(n8148), .B2(n5889), .ZN(n6173)
         );
  OAI221_X1 U4127 ( .B1(n897), .B2(n5890), .C1(n961), .C2(n5891), .A(n6174), 
        .ZN(n6167) );
  AOI222_X1 U4128 ( .A1(n5893), .A2(n4927), .B1(n5894), .B2(n5186), .C1(n5895), 
        .C2(n5525), .ZN(n6174) );
  OAI22_X1 U4129 ( .A1(n7893), .A2(n5870), .B1(n6175), .B2(n5872), .ZN(n8343)
         );
  NOR4_X1 U4130 ( .A1(n6176), .A2(n6177), .A3(n6178), .A4(n6179), .ZN(n6175)
         );
  OAI221_X1 U4131 ( .B1(n5830), .B2(n4862), .C1(n5877), .C2(n5057), .A(n6180), 
        .ZN(n6179) );
  AOI22_X1 U4132 ( .A1(n5879), .A2(n5267), .B1(n5880), .B2(n4992), .ZN(n6180)
         );
  OAI221_X1 U4133 ( .B1(n514), .B2(n5881), .C1(n578), .C2(n5882), .A(n6181), 
        .ZN(n6178) );
  AOI22_X1 U4134 ( .A1(n8085), .A2(n5884), .B1(n8021), .B2(n5885), .ZN(n6181)
         );
  OAI221_X1 U4135 ( .B1(n770), .B2(n5819), .C1(n834), .C2(n5886), .A(n6182), 
        .ZN(n6177) );
  AOI22_X1 U4136 ( .A1(n8213), .A2(n5888), .B1(n8149), .B2(n5889), .ZN(n6182)
         );
  OAI221_X1 U4137 ( .B1(n898), .B2(n5890), .C1(n962), .C2(n5891), .A(n6183), 
        .ZN(n6176) );
  AOI222_X1 U4138 ( .A1(n5893), .A2(n4926), .B1(n5894), .B2(n5185), .C1(n5895), 
        .C2(n5524), .ZN(n6183) );
  OAI22_X1 U4139 ( .A1(n7894), .A2(n5870), .B1(n6184), .B2(n5872), .ZN(n8344)
         );
  NOR4_X1 U4140 ( .A1(n6185), .A2(n6186), .A3(n6187), .A4(n6188), .ZN(n6184)
         );
  OAI221_X1 U4141 ( .B1(n5830), .B2(n4861), .C1(n5877), .C2(n5056), .A(n6189), 
        .ZN(n6188) );
  AOI22_X1 U4142 ( .A1(n5879), .A2(n5266), .B1(n5880), .B2(n4991), .ZN(n6189)
         );
  OAI221_X1 U4143 ( .B1(n515), .B2(n5881), .C1(n579), .C2(n5882), .A(n6190), 
        .ZN(n6187) );
  AOI22_X1 U4144 ( .A1(n8086), .A2(n5884), .B1(n8022), .B2(n5885), .ZN(n6190)
         );
  OAI221_X1 U4145 ( .B1(n771), .B2(n5819), .C1(n835), .C2(n5886), .A(n6191), 
        .ZN(n6186) );
  AOI22_X1 U4146 ( .A1(n8214), .A2(n5888), .B1(n8150), .B2(n5889), .ZN(n6191)
         );
  OAI221_X1 U4147 ( .B1(n899), .B2(n5890), .C1(n963), .C2(n5891), .A(n6192), 
        .ZN(n6185) );
  AOI222_X1 U4148 ( .A1(n5893), .A2(n4925), .B1(n5894), .B2(n5184), .C1(n5895), 
        .C2(n5523), .ZN(n6192) );
  OAI22_X1 U4149 ( .A1(n7895), .A2(n5870), .B1(n6193), .B2(n5872), .ZN(n8345)
         );
  NOR4_X1 U4150 ( .A1(n6194), .A2(n6195), .A3(n6196), .A4(n6197), .ZN(n6193)
         );
  OAI221_X1 U4151 ( .B1(n5830), .B2(n4860), .C1(n5877), .C2(n5055), .A(n6198), 
        .ZN(n6197) );
  AOI22_X1 U4152 ( .A1(n5879), .A2(n5265), .B1(n5880), .B2(n4990), .ZN(n6198)
         );
  OAI221_X1 U4153 ( .B1(n516), .B2(n5881), .C1(n580), .C2(n5882), .A(n6199), 
        .ZN(n6196) );
  AOI22_X1 U4154 ( .A1(n8087), .A2(n5884), .B1(n8023), .B2(n5885), .ZN(n6199)
         );
  OAI221_X1 U4155 ( .B1(n772), .B2(n5819), .C1(n836), .C2(n5886), .A(n6200), 
        .ZN(n6195) );
  AOI22_X1 U4156 ( .A1(n8215), .A2(n5888), .B1(n8151), .B2(n5889), .ZN(n6200)
         );
  OAI221_X1 U4157 ( .B1(n900), .B2(n5890), .C1(n964), .C2(n5891), .A(n6201), 
        .ZN(n6194) );
  AOI222_X1 U4158 ( .A1(n5893), .A2(n4924), .B1(n5894), .B2(n5183), .C1(n5895), 
        .C2(n5522), .ZN(n6201) );
  OAI22_X1 U4159 ( .A1(n7896), .A2(n5870), .B1(n6202), .B2(n5872), .ZN(n8346)
         );
  NOR4_X1 U4160 ( .A1(n6203), .A2(n6204), .A3(n6205), .A4(n6206), .ZN(n6202)
         );
  OAI221_X1 U4161 ( .B1(n5830), .B2(n4859), .C1(n5877), .C2(n5054), .A(n6207), 
        .ZN(n6206) );
  AOI22_X1 U4162 ( .A1(n5879), .A2(n5264), .B1(n5880), .B2(n4989), .ZN(n6207)
         );
  OAI221_X1 U4163 ( .B1(n517), .B2(n5881), .C1(n581), .C2(n5882), .A(n6208), 
        .ZN(n6205) );
  AOI22_X1 U4164 ( .A1(n8088), .A2(n5884), .B1(n8024), .B2(n5885), .ZN(n6208)
         );
  OAI221_X1 U4165 ( .B1(n773), .B2(n5819), .C1(n837), .C2(n5886), .A(n6209), 
        .ZN(n6204) );
  AOI22_X1 U4166 ( .A1(n8216), .A2(n5888), .B1(n8152), .B2(n5889), .ZN(n6209)
         );
  OAI221_X1 U4167 ( .B1(n901), .B2(n5890), .C1(n965), .C2(n5891), .A(n6210), 
        .ZN(n6203) );
  AOI222_X1 U4168 ( .A1(n5893), .A2(n4923), .B1(n5894), .B2(n5182), .C1(n5895), 
        .C2(n5521), .ZN(n6210) );
  OAI22_X1 U4169 ( .A1(n7897), .A2(n5870), .B1(n6211), .B2(n5872), .ZN(n8347)
         );
  NOR4_X1 U4170 ( .A1(n6212), .A2(n6213), .A3(n6214), .A4(n6215), .ZN(n6211)
         );
  OAI221_X1 U4171 ( .B1(n5830), .B2(n4858), .C1(n5877), .C2(n5053), .A(n6216), 
        .ZN(n6215) );
  AOI22_X1 U4172 ( .A1(n5879), .A2(n5263), .B1(n5880), .B2(n4988), .ZN(n6216)
         );
  OAI221_X1 U4173 ( .B1(n518), .B2(n5881), .C1(n582), .C2(n5882), .A(n6217), 
        .ZN(n6214) );
  AOI22_X1 U4174 ( .A1(n8089), .A2(n5884), .B1(n8025), .B2(n5885), .ZN(n6217)
         );
  OAI221_X1 U4175 ( .B1(n774), .B2(n5819), .C1(n838), .C2(n5886), .A(n6218), 
        .ZN(n6213) );
  AOI22_X1 U4176 ( .A1(n8217), .A2(n5888), .B1(n8153), .B2(n5889), .ZN(n6218)
         );
  OAI221_X1 U4177 ( .B1(n902), .B2(n5890), .C1(n966), .C2(n5891), .A(n6219), 
        .ZN(n6212) );
  AOI222_X1 U4178 ( .A1(n5893), .A2(n4922), .B1(n5894), .B2(n5181), .C1(n5895), 
        .C2(n5520), .ZN(n6219) );
  OAI22_X1 U4179 ( .A1(n7898), .A2(n5870), .B1(n6220), .B2(n5872), .ZN(n8348)
         );
  NOR4_X1 U4180 ( .A1(n6221), .A2(n6222), .A3(n6223), .A4(n6224), .ZN(n6220)
         );
  OAI221_X1 U4181 ( .B1(n5830), .B2(n4857), .C1(n5877), .C2(n5052), .A(n6225), 
        .ZN(n6224) );
  AOI22_X1 U4182 ( .A1(n5879), .A2(n5262), .B1(n5880), .B2(n4987), .ZN(n6225)
         );
  OAI221_X1 U4183 ( .B1(n519), .B2(n5881), .C1(n583), .C2(n5882), .A(n6226), 
        .ZN(n6223) );
  AOI22_X1 U4184 ( .A1(n8090), .A2(n5884), .B1(n8026), .B2(n5885), .ZN(n6226)
         );
  OAI221_X1 U4185 ( .B1(n775), .B2(n5819), .C1(n839), .C2(n5886), .A(n6227), 
        .ZN(n6222) );
  AOI22_X1 U4186 ( .A1(n8218), .A2(n5888), .B1(n8154), .B2(n5889), .ZN(n6227)
         );
  OAI221_X1 U4187 ( .B1(n903), .B2(n5890), .C1(n967), .C2(n5891), .A(n6228), 
        .ZN(n6221) );
  AOI222_X1 U4188 ( .A1(n5893), .A2(n4921), .B1(n5894), .B2(n5180), .C1(n5895), 
        .C2(n5519), .ZN(n6228) );
  OAI22_X1 U4189 ( .A1(n7899), .A2(n5870), .B1(n6229), .B2(n5872), .ZN(n8349)
         );
  NOR4_X1 U4190 ( .A1(n6230), .A2(n6231), .A3(n6232), .A4(n6233), .ZN(n6229)
         );
  OAI221_X1 U4191 ( .B1(n5830), .B2(n4856), .C1(n5877), .C2(n5051), .A(n6234), 
        .ZN(n6233) );
  AOI22_X1 U4192 ( .A1(n5879), .A2(n5261), .B1(n5880), .B2(n4986), .ZN(n6234)
         );
  OAI221_X1 U4193 ( .B1(n520), .B2(n5881), .C1(n584), .C2(n5882), .A(n6235), 
        .ZN(n6232) );
  AOI22_X1 U4194 ( .A1(n8091), .A2(n5884), .B1(n8027), .B2(n5885), .ZN(n6235)
         );
  OAI221_X1 U4195 ( .B1(n776), .B2(n5819), .C1(n840), .C2(n5886), .A(n6236), 
        .ZN(n6231) );
  AOI22_X1 U4196 ( .A1(n8219), .A2(n5888), .B1(n8155), .B2(n5889), .ZN(n6236)
         );
  OAI221_X1 U4197 ( .B1(n904), .B2(n5890), .C1(n968), .C2(n5891), .A(n6237), 
        .ZN(n6230) );
  AOI222_X1 U4198 ( .A1(n5893), .A2(n4920), .B1(n5894), .B2(n5179), .C1(n5895), 
        .C2(n5518), .ZN(n6237) );
  OAI22_X1 U4199 ( .A1(n7900), .A2(n5870), .B1(n6238), .B2(n5872), .ZN(n8350)
         );
  NOR4_X1 U4200 ( .A1(n6239), .A2(n6240), .A3(n6241), .A4(n6242), .ZN(n6238)
         );
  OAI221_X1 U4201 ( .B1(n5830), .B2(n4855), .C1(n5877), .C2(n5050), .A(n6243), 
        .ZN(n6242) );
  AOI22_X1 U4202 ( .A1(n5879), .A2(n5260), .B1(n5880), .B2(n4985), .ZN(n6243)
         );
  OAI221_X1 U4203 ( .B1(n521), .B2(n5881), .C1(n585), .C2(n5882), .A(n6244), 
        .ZN(n6241) );
  AOI22_X1 U4204 ( .A1(n8092), .A2(n5884), .B1(n8028), .B2(n5885), .ZN(n6244)
         );
  OAI221_X1 U4205 ( .B1(n777), .B2(n5819), .C1(n841), .C2(n5886), .A(n6245), 
        .ZN(n6240) );
  AOI22_X1 U4206 ( .A1(n8220), .A2(n5888), .B1(n8156), .B2(n5889), .ZN(n6245)
         );
  OAI221_X1 U4207 ( .B1(n905), .B2(n5890), .C1(n969), .C2(n5891), .A(n6246), 
        .ZN(n6239) );
  AOI222_X1 U4208 ( .A1(n5893), .A2(n4919), .B1(n5894), .B2(n5178), .C1(n5895), 
        .C2(n5517), .ZN(n6246) );
  OAI22_X1 U4209 ( .A1(n7901), .A2(n5870), .B1(n6247), .B2(n5872), .ZN(n8351)
         );
  NOR4_X1 U4210 ( .A1(n6248), .A2(n6249), .A3(n6250), .A4(n6251), .ZN(n6247)
         );
  OAI221_X1 U4211 ( .B1(n5830), .B2(n4854), .C1(n5877), .C2(n5049), .A(n6252), 
        .ZN(n6251) );
  AOI22_X1 U4212 ( .A1(n5879), .A2(n5259), .B1(n5880), .B2(n4984), .ZN(n6252)
         );
  OAI221_X1 U4213 ( .B1(n522), .B2(n5881), .C1(n586), .C2(n5882), .A(n6253), 
        .ZN(n6250) );
  AOI22_X1 U4214 ( .A1(n8093), .A2(n5884), .B1(n8029), .B2(n5885), .ZN(n6253)
         );
  OAI221_X1 U4215 ( .B1(n778), .B2(n5819), .C1(n842), .C2(n5886), .A(n6254), 
        .ZN(n6249) );
  AOI22_X1 U4216 ( .A1(n8221), .A2(n5888), .B1(n8157), .B2(n5889), .ZN(n6254)
         );
  OAI221_X1 U4217 ( .B1(n906), .B2(n5890), .C1(n970), .C2(n5891), .A(n6255), 
        .ZN(n6248) );
  AOI222_X1 U4218 ( .A1(n5893), .A2(n4918), .B1(n5894), .B2(n5177), .C1(n5895), 
        .C2(n5516), .ZN(n6255) );
  OAI22_X1 U4219 ( .A1(n7902), .A2(n5870), .B1(n6256), .B2(n5872), .ZN(n8352)
         );
  NOR4_X1 U4220 ( .A1(n6257), .A2(n6258), .A3(n6259), .A4(n6260), .ZN(n6256)
         );
  OAI221_X1 U4221 ( .B1(n5830), .B2(n4853), .C1(n5877), .C2(n5048), .A(n6261), 
        .ZN(n6260) );
  AOI22_X1 U4222 ( .A1(n5879), .A2(n5258), .B1(n5880), .B2(n4983), .ZN(n6261)
         );
  OAI221_X1 U4223 ( .B1(n523), .B2(n5881), .C1(n587), .C2(n5882), .A(n6262), 
        .ZN(n6259) );
  AOI22_X1 U4224 ( .A1(n8094), .A2(n5884), .B1(n8030), .B2(n5885), .ZN(n6262)
         );
  OAI221_X1 U4225 ( .B1(n779), .B2(n5819), .C1(n843), .C2(n5886), .A(n6263), 
        .ZN(n6258) );
  AOI22_X1 U4226 ( .A1(n8222), .A2(n5888), .B1(n8158), .B2(n5889), .ZN(n6263)
         );
  OAI221_X1 U4227 ( .B1(n907), .B2(n5890), .C1(n971), .C2(n5891), .A(n6264), 
        .ZN(n6257) );
  AOI222_X1 U4228 ( .A1(n5893), .A2(n4917), .B1(n5894), .B2(n5176), .C1(n5895), 
        .C2(n5515), .ZN(n6264) );
  OAI22_X1 U4229 ( .A1(n7903), .A2(n5870), .B1(n6265), .B2(n5872), .ZN(n8353)
         );
  NOR4_X1 U4230 ( .A1(n6266), .A2(n6267), .A3(n6268), .A4(n6269), .ZN(n6265)
         );
  OAI221_X1 U4231 ( .B1(n5830), .B2(n4852), .C1(n5877), .C2(n5047), .A(n6270), 
        .ZN(n6269) );
  AOI22_X1 U4232 ( .A1(n5879), .A2(n5257), .B1(n5880), .B2(n4982), .ZN(n6270)
         );
  OAI221_X1 U4233 ( .B1(n524), .B2(n5881), .C1(n588), .C2(n5882), .A(n6271), 
        .ZN(n6268) );
  AOI22_X1 U4234 ( .A1(n8095), .A2(n5884), .B1(n8031), .B2(n5885), .ZN(n6271)
         );
  OAI221_X1 U4235 ( .B1(n780), .B2(n5819), .C1(n844), .C2(n5886), .A(n6272), 
        .ZN(n6267) );
  AOI22_X1 U4236 ( .A1(n8223), .A2(n5888), .B1(n8159), .B2(n5889), .ZN(n6272)
         );
  OAI221_X1 U4237 ( .B1(n908), .B2(n5890), .C1(n972), .C2(n5891), .A(n6273), 
        .ZN(n6266) );
  AOI222_X1 U4238 ( .A1(n5893), .A2(n4916), .B1(n5894), .B2(n5175), .C1(n5895), 
        .C2(n5514), .ZN(n6273) );
  OAI22_X1 U4239 ( .A1(n7904), .A2(n5870), .B1(n6274), .B2(n5872), .ZN(n8354)
         );
  NOR4_X1 U4240 ( .A1(n6275), .A2(n6276), .A3(n6277), .A4(n6278), .ZN(n6274)
         );
  OAI221_X1 U4241 ( .B1(n5830), .B2(n4851), .C1(n5877), .C2(n5046), .A(n6279), 
        .ZN(n6278) );
  AOI22_X1 U4242 ( .A1(n5879), .A2(n5256), .B1(n5880), .B2(n4981), .ZN(n6279)
         );
  OAI221_X1 U4243 ( .B1(n525), .B2(n5881), .C1(n589), .C2(n5882), .A(n6280), 
        .ZN(n6277) );
  AOI22_X1 U4244 ( .A1(n8096), .A2(n5884), .B1(n8032), .B2(n5885), .ZN(n6280)
         );
  OAI221_X1 U4245 ( .B1(n781), .B2(n5819), .C1(n845), .C2(n5886), .A(n6281), 
        .ZN(n6276) );
  AOI22_X1 U4246 ( .A1(n8224), .A2(n5888), .B1(n8160), .B2(n5889), .ZN(n6281)
         );
  OAI221_X1 U4247 ( .B1(n909), .B2(n5890), .C1(n973), .C2(n5891), .A(n6282), 
        .ZN(n6275) );
  AOI222_X1 U4248 ( .A1(n5893), .A2(n4915), .B1(n5894), .B2(n5174), .C1(n5895), 
        .C2(n5513), .ZN(n6282) );
  OAI22_X1 U4249 ( .A1(n7905), .A2(n5870), .B1(n6283), .B2(n5872), .ZN(n8355)
         );
  NOR4_X1 U4250 ( .A1(n6284), .A2(n6285), .A3(n6286), .A4(n6287), .ZN(n6283)
         );
  OAI221_X1 U4251 ( .B1(n5830), .B2(n4850), .C1(n5877), .C2(n5045), .A(n6288), 
        .ZN(n6287) );
  AOI22_X1 U4252 ( .A1(n5879), .A2(n5255), .B1(n5880), .B2(n4980), .ZN(n6288)
         );
  OAI221_X1 U4253 ( .B1(n526), .B2(n5881), .C1(n590), .C2(n5882), .A(n6289), 
        .ZN(n6286) );
  AOI22_X1 U4254 ( .A1(n8097), .A2(n5884), .B1(n8033), .B2(n5885), .ZN(n6289)
         );
  OAI221_X1 U4255 ( .B1(n782), .B2(n5819), .C1(n846), .C2(n5886), .A(n6290), 
        .ZN(n6285) );
  AOI22_X1 U4256 ( .A1(n8225), .A2(n5888), .B1(n8161), .B2(n5889), .ZN(n6290)
         );
  OAI221_X1 U4257 ( .B1(n910), .B2(n5890), .C1(n974), .C2(n5891), .A(n6291), 
        .ZN(n6284) );
  AOI222_X1 U4258 ( .A1(n5893), .A2(n4914), .B1(n5894), .B2(n5173), .C1(n5895), 
        .C2(n5512), .ZN(n6291) );
  OAI22_X1 U4259 ( .A1(n7906), .A2(n5870), .B1(n6292), .B2(n5872), .ZN(n8356)
         );
  NOR4_X1 U4260 ( .A1(n6293), .A2(n6294), .A3(n6295), .A4(n6296), .ZN(n6292)
         );
  OAI221_X1 U4261 ( .B1(n5830), .B2(n4849), .C1(n5877), .C2(n5044), .A(n6297), 
        .ZN(n6296) );
  AOI22_X1 U4262 ( .A1(n5879), .A2(n5254), .B1(n5880), .B2(n4979), .ZN(n6297)
         );
  OAI221_X1 U4263 ( .B1(n527), .B2(n5881), .C1(n591), .C2(n5882), .A(n6298), 
        .ZN(n6295) );
  AOI22_X1 U4264 ( .A1(n8098), .A2(n5884), .B1(n8034), .B2(n5885), .ZN(n6298)
         );
  OAI221_X1 U4265 ( .B1(n783), .B2(n5819), .C1(n847), .C2(n5886), .A(n6299), 
        .ZN(n6294) );
  AOI22_X1 U4266 ( .A1(n8226), .A2(n5888), .B1(n8162), .B2(n5889), .ZN(n6299)
         );
  OAI221_X1 U4267 ( .B1(n911), .B2(n5890), .C1(n975), .C2(n5891), .A(n6300), 
        .ZN(n6293) );
  AOI222_X1 U4268 ( .A1(n5893), .A2(n4913), .B1(n5894), .B2(n5172), .C1(n5895), 
        .C2(n5511), .ZN(n6300) );
  OAI22_X1 U4269 ( .A1(n7907), .A2(n5870), .B1(n6301), .B2(n5872), .ZN(n8357)
         );
  NOR4_X1 U4270 ( .A1(n6302), .A2(n6303), .A3(n6304), .A4(n6305), .ZN(n6301)
         );
  OAI221_X1 U4271 ( .B1(n5830), .B2(n4848), .C1(n5877), .C2(n5043), .A(n6306), 
        .ZN(n6305) );
  AOI22_X1 U4272 ( .A1(n5879), .A2(n5253), .B1(n5880), .B2(n4978), .ZN(n6306)
         );
  OAI221_X1 U4273 ( .B1(n528), .B2(n5881), .C1(n592), .C2(n5882), .A(n6307), 
        .ZN(n6304) );
  AOI22_X1 U4274 ( .A1(n8099), .A2(n5884), .B1(n8035), .B2(n5885), .ZN(n6307)
         );
  OAI221_X1 U4275 ( .B1(n784), .B2(n5819), .C1(n848), .C2(n5886), .A(n6308), 
        .ZN(n6303) );
  AOI22_X1 U4276 ( .A1(n8227), .A2(n5888), .B1(n8163), .B2(n5889), .ZN(n6308)
         );
  OAI221_X1 U4277 ( .B1(n912), .B2(n5890), .C1(n976), .C2(n5891), .A(n6309), 
        .ZN(n6302) );
  AOI222_X1 U4278 ( .A1(n5893), .A2(n4912), .B1(n5894), .B2(n5171), .C1(n5895), 
        .C2(n5510), .ZN(n6309) );
  OAI22_X1 U4279 ( .A1(n7908), .A2(n5870), .B1(n6310), .B2(n5872), .ZN(n8358)
         );
  NOR4_X1 U4280 ( .A1(n6311), .A2(n6312), .A3(n6313), .A4(n6314), .ZN(n6310)
         );
  OAI221_X1 U4281 ( .B1(n5830), .B2(n4847), .C1(n5877), .C2(n5042), .A(n6315), 
        .ZN(n6314) );
  AOI22_X1 U4282 ( .A1(n5879), .A2(n5252), .B1(n5880), .B2(n4977), .ZN(n6315)
         );
  OAI221_X1 U4283 ( .B1(n529), .B2(n5881), .C1(n593), .C2(n5882), .A(n6316), 
        .ZN(n6313) );
  AOI22_X1 U4284 ( .A1(n8100), .A2(n5884), .B1(n8036), .B2(n5885), .ZN(n6316)
         );
  OAI221_X1 U4285 ( .B1(n785), .B2(n5819), .C1(n849), .C2(n5886), .A(n6317), 
        .ZN(n6312) );
  AOI22_X1 U4286 ( .A1(n8228), .A2(n5888), .B1(n8164), .B2(n5889), .ZN(n6317)
         );
  OAI221_X1 U4287 ( .B1(n913), .B2(n5890), .C1(n977), .C2(n5891), .A(n6318), 
        .ZN(n6311) );
  AOI222_X1 U4288 ( .A1(n5893), .A2(n4911), .B1(n5894), .B2(n5170), .C1(n5895), 
        .C2(n5509), .ZN(n6318) );
  OAI22_X1 U4289 ( .A1(n7909), .A2(n5870), .B1(n6319), .B2(n5872), .ZN(n8359)
         );
  NOR4_X1 U4290 ( .A1(n6320), .A2(n6321), .A3(n6322), .A4(n6323), .ZN(n6319)
         );
  OAI221_X1 U4291 ( .B1(n5830), .B2(n4846), .C1(n5877), .C2(n5041), .A(n6324), 
        .ZN(n6323) );
  AOI22_X1 U4292 ( .A1(n5879), .A2(n5251), .B1(n5880), .B2(n4976), .ZN(n6324)
         );
  OAI221_X1 U4293 ( .B1(n530), .B2(n5881), .C1(n594), .C2(n5882), .A(n6325), 
        .ZN(n6322) );
  AOI22_X1 U4294 ( .A1(n8101), .A2(n5884), .B1(n8037), .B2(n5885), .ZN(n6325)
         );
  OAI221_X1 U4295 ( .B1(n786), .B2(n5819), .C1(n850), .C2(n5886), .A(n6326), 
        .ZN(n6321) );
  AOI22_X1 U4296 ( .A1(n8229), .A2(n5888), .B1(n8165), .B2(n5889), .ZN(n6326)
         );
  OAI221_X1 U4297 ( .B1(n914), .B2(n5890), .C1(n978), .C2(n5891), .A(n6327), 
        .ZN(n6320) );
  AOI222_X1 U4298 ( .A1(n5893), .A2(n4910), .B1(n5894), .B2(n5169), .C1(n5895), 
        .C2(n5508), .ZN(n6327) );
  OAI22_X1 U4299 ( .A1(n7910), .A2(n5870), .B1(n6328), .B2(n5872), .ZN(n8360)
         );
  NOR4_X1 U4300 ( .A1(n6329), .A2(n6330), .A3(n6331), .A4(n6332), .ZN(n6328)
         );
  OAI221_X1 U4301 ( .B1(n5830), .B2(n4845), .C1(n5877), .C2(n5040), .A(n6333), 
        .ZN(n6332) );
  AOI22_X1 U4302 ( .A1(n5879), .A2(n5250), .B1(n5880), .B2(n4975), .ZN(n6333)
         );
  OAI221_X1 U4303 ( .B1(n531), .B2(n5881), .C1(n595), .C2(n5882), .A(n6334), 
        .ZN(n6331) );
  AOI22_X1 U4304 ( .A1(n8102), .A2(n5884), .B1(n8038), .B2(n5885), .ZN(n6334)
         );
  OAI221_X1 U4305 ( .B1(n787), .B2(n5819), .C1(n851), .C2(n5886), .A(n6335), 
        .ZN(n6330) );
  AOI22_X1 U4306 ( .A1(n8230), .A2(n5888), .B1(n8166), .B2(n5889), .ZN(n6335)
         );
  OAI221_X1 U4307 ( .B1(n915), .B2(n5890), .C1(n979), .C2(n5891), .A(n6336), 
        .ZN(n6329) );
  AOI222_X1 U4308 ( .A1(n5893), .A2(n4909), .B1(n5894), .B2(n5168), .C1(n5895), 
        .C2(n5507), .ZN(n6336) );
  OAI22_X1 U4309 ( .A1(n7911), .A2(n5870), .B1(n6337), .B2(n5872), .ZN(n8361)
         );
  NOR4_X1 U4310 ( .A1(n6338), .A2(n6339), .A3(n6340), .A4(n6341), .ZN(n6337)
         );
  OAI221_X1 U4311 ( .B1(n5830), .B2(n4844), .C1(n5877), .C2(n5039), .A(n6342), 
        .ZN(n6341) );
  AOI22_X1 U4312 ( .A1(n5879), .A2(n5249), .B1(n5880), .B2(n4974), .ZN(n6342)
         );
  OAI221_X1 U4313 ( .B1(n532), .B2(n5881), .C1(n596), .C2(n5882), .A(n6343), 
        .ZN(n6340) );
  AOI22_X1 U4314 ( .A1(n8103), .A2(n5884), .B1(n8039), .B2(n5885), .ZN(n6343)
         );
  OAI221_X1 U4315 ( .B1(n788), .B2(n5819), .C1(n852), .C2(n5886), .A(n6344), 
        .ZN(n6339) );
  AOI22_X1 U4316 ( .A1(n8231), .A2(n5888), .B1(n8167), .B2(n5889), .ZN(n6344)
         );
  OAI221_X1 U4317 ( .B1(n916), .B2(n5890), .C1(n980), .C2(n5891), .A(n6345), 
        .ZN(n6338) );
  AOI222_X1 U4318 ( .A1(n5893), .A2(n4908), .B1(n5894), .B2(n5167), .C1(n5895), 
        .C2(n5506), .ZN(n6345) );
  OAI22_X1 U4319 ( .A1(n7912), .A2(n5870), .B1(n6346), .B2(n5872), .ZN(n8362)
         );
  NOR4_X1 U4320 ( .A1(n6347), .A2(n6348), .A3(n6349), .A4(n6350), .ZN(n6346)
         );
  OAI221_X1 U4321 ( .B1(n5830), .B2(n4843), .C1(n5877), .C2(n5038), .A(n6351), 
        .ZN(n6350) );
  AOI22_X1 U4322 ( .A1(n5879), .A2(n5248), .B1(n5880), .B2(n4973), .ZN(n6351)
         );
  OAI221_X1 U4323 ( .B1(n533), .B2(n5881), .C1(n597), .C2(n5882), .A(n6352), 
        .ZN(n6349) );
  AOI22_X1 U4324 ( .A1(n8104), .A2(n5884), .B1(n8040), .B2(n5885), .ZN(n6352)
         );
  OAI221_X1 U4325 ( .B1(n789), .B2(n5819), .C1(n853), .C2(n5886), .A(n6353), 
        .ZN(n6348) );
  AOI22_X1 U4326 ( .A1(n8232), .A2(n5888), .B1(n8168), .B2(n5889), .ZN(n6353)
         );
  OAI221_X1 U4327 ( .B1(n917), .B2(n5890), .C1(n981), .C2(n5891), .A(n6354), 
        .ZN(n6347) );
  AOI222_X1 U4328 ( .A1(n5893), .A2(n4907), .B1(n5894), .B2(n5166), .C1(n5895), 
        .C2(n5505), .ZN(n6354) );
  OAI22_X1 U4329 ( .A1(n7913), .A2(n5870), .B1(n6355), .B2(n5872), .ZN(n8363)
         );
  NOR4_X1 U4330 ( .A1(n6356), .A2(n6357), .A3(n6358), .A4(n6359), .ZN(n6355)
         );
  OAI221_X1 U4331 ( .B1(n5830), .B2(n4842), .C1(n5877), .C2(n5037), .A(n6360), 
        .ZN(n6359) );
  AOI22_X1 U4332 ( .A1(n5879), .A2(n5247), .B1(n5880), .B2(n4972), .ZN(n6360)
         );
  OAI221_X1 U4333 ( .B1(n534), .B2(n5881), .C1(n598), .C2(n5882), .A(n6361), 
        .ZN(n6358) );
  AOI22_X1 U4334 ( .A1(n8105), .A2(n5884), .B1(n8041), .B2(n5885), .ZN(n6361)
         );
  OAI221_X1 U4335 ( .B1(n790), .B2(n5819), .C1(n854), .C2(n5886), .A(n6362), 
        .ZN(n6357) );
  AOI22_X1 U4336 ( .A1(n8233), .A2(n5888), .B1(n8169), .B2(n5889), .ZN(n6362)
         );
  OAI221_X1 U4337 ( .B1(n918), .B2(n5890), .C1(n982), .C2(n5891), .A(n6363), 
        .ZN(n6356) );
  AOI222_X1 U4338 ( .A1(n5893), .A2(n4906), .B1(n5894), .B2(n5165), .C1(n5895), 
        .C2(n5504), .ZN(n6363) );
  OAI22_X1 U4339 ( .A1(n7914), .A2(n5870), .B1(n6364), .B2(n5872), .ZN(n8364)
         );
  NOR4_X1 U4340 ( .A1(n6365), .A2(n6366), .A3(n6367), .A4(n6368), .ZN(n6364)
         );
  OAI221_X1 U4341 ( .B1(n5830), .B2(n4841), .C1(n5877), .C2(n5036), .A(n6369), 
        .ZN(n6368) );
  AOI22_X1 U4342 ( .A1(n5879), .A2(n5246), .B1(n5880), .B2(n4971), .ZN(n6369)
         );
  OAI221_X1 U4343 ( .B1(n535), .B2(n5881), .C1(n599), .C2(n5882), .A(n6370), 
        .ZN(n6367) );
  AOI22_X1 U4344 ( .A1(n8106), .A2(n5884), .B1(n8042), .B2(n5885), .ZN(n6370)
         );
  OAI221_X1 U4345 ( .B1(n791), .B2(n5819), .C1(n855), .C2(n5886), .A(n6371), 
        .ZN(n6366) );
  AOI22_X1 U4346 ( .A1(n8234), .A2(n5888), .B1(n8170), .B2(n5889), .ZN(n6371)
         );
  OAI221_X1 U4347 ( .B1(n919), .B2(n5890), .C1(n983), .C2(n5891), .A(n6372), 
        .ZN(n6365) );
  AOI222_X1 U4348 ( .A1(n5893), .A2(n4905), .B1(n5894), .B2(n5164), .C1(n5895), 
        .C2(n5503), .ZN(n6372) );
  OAI22_X1 U4349 ( .A1(n7915), .A2(n5870), .B1(n6373), .B2(n5872), .ZN(n8365)
         );
  NOR4_X1 U4350 ( .A1(n6374), .A2(n6375), .A3(n6376), .A4(n6377), .ZN(n6373)
         );
  OAI221_X1 U4351 ( .B1(n5830), .B2(n4840), .C1(n5877), .C2(n5035), .A(n6378), 
        .ZN(n6377) );
  AOI22_X1 U4352 ( .A1(n5879), .A2(n5245), .B1(n5880), .B2(n4970), .ZN(n6378)
         );
  OAI221_X1 U4353 ( .B1(n536), .B2(n5881), .C1(n600), .C2(n5882), .A(n6379), 
        .ZN(n6376) );
  AOI22_X1 U4354 ( .A1(n8107), .A2(n5884), .B1(n8043), .B2(n5885), .ZN(n6379)
         );
  OAI221_X1 U4355 ( .B1(n792), .B2(n5819), .C1(n856), .C2(n5886), .A(n6380), 
        .ZN(n6375) );
  AOI22_X1 U4356 ( .A1(n8235), .A2(n5888), .B1(n8171), .B2(n5889), .ZN(n6380)
         );
  OAI221_X1 U4357 ( .B1(n920), .B2(n5890), .C1(n984), .C2(n5891), .A(n6381), 
        .ZN(n6374) );
  AOI222_X1 U4358 ( .A1(n5893), .A2(n4904), .B1(n5894), .B2(n5163), .C1(n5895), 
        .C2(n5502), .ZN(n6381) );
  OAI22_X1 U4359 ( .A1(n7916), .A2(n5870), .B1(n6382), .B2(n5872), .ZN(n8366)
         );
  NOR4_X1 U4360 ( .A1(n6383), .A2(n6384), .A3(n6385), .A4(n6386), .ZN(n6382)
         );
  OAI221_X1 U4361 ( .B1(n5830), .B2(n4839), .C1(n5877), .C2(n5034), .A(n6387), 
        .ZN(n6386) );
  AOI22_X1 U4362 ( .A1(n5879), .A2(n5244), .B1(n5880), .B2(n4969), .ZN(n6387)
         );
  OAI221_X1 U4363 ( .B1(n537), .B2(n5881), .C1(n601), .C2(n5882), .A(n6388), 
        .ZN(n6385) );
  AOI22_X1 U4364 ( .A1(n8108), .A2(n5884), .B1(n8044), .B2(n5885), .ZN(n6388)
         );
  OAI221_X1 U4365 ( .B1(n793), .B2(n5819), .C1(n857), .C2(n5886), .A(n6389), 
        .ZN(n6384) );
  AOI22_X1 U4366 ( .A1(n8236), .A2(n5888), .B1(n8172), .B2(n5889), .ZN(n6389)
         );
  OAI221_X1 U4367 ( .B1(n921), .B2(n5890), .C1(n985), .C2(n5891), .A(n6390), 
        .ZN(n6383) );
  AOI222_X1 U4368 ( .A1(n5893), .A2(n4903), .B1(n5894), .B2(n5162), .C1(n5895), 
        .C2(n5501), .ZN(n6390) );
  OAI22_X1 U4369 ( .A1(n7917), .A2(n5870), .B1(n6391), .B2(n5872), .ZN(n8367)
         );
  NOR4_X1 U4370 ( .A1(n6392), .A2(n6393), .A3(n6394), .A4(n6395), .ZN(n6391)
         );
  OAI221_X1 U4371 ( .B1(n5830), .B2(n4838), .C1(n5877), .C2(n5033), .A(n6396), 
        .ZN(n6395) );
  AOI22_X1 U4372 ( .A1(n5879), .A2(n5243), .B1(n5880), .B2(n4968), .ZN(n6396)
         );
  OAI221_X1 U4373 ( .B1(n538), .B2(n5881), .C1(n602), .C2(n5882), .A(n6397), 
        .ZN(n6394) );
  AOI22_X1 U4374 ( .A1(n8109), .A2(n5884), .B1(n8045), .B2(n5885), .ZN(n6397)
         );
  OAI221_X1 U4375 ( .B1(n794), .B2(n5819), .C1(n858), .C2(n5886), .A(n6398), 
        .ZN(n6393) );
  AOI22_X1 U4376 ( .A1(n8237), .A2(n5888), .B1(n8173), .B2(n5889), .ZN(n6398)
         );
  OAI221_X1 U4377 ( .B1(n922), .B2(n5890), .C1(n986), .C2(n5891), .A(n6399), 
        .ZN(n6392) );
  AOI222_X1 U4378 ( .A1(n5893), .A2(n4902), .B1(n5894), .B2(n5161), .C1(n5895), 
        .C2(n5500), .ZN(n6399) );
  OAI22_X1 U4379 ( .A1(n7918), .A2(n5870), .B1(n6400), .B2(n5872), .ZN(n8368)
         );
  NOR4_X1 U4380 ( .A1(n6401), .A2(n6402), .A3(n6403), .A4(n6404), .ZN(n6400)
         );
  OAI221_X1 U4381 ( .B1(n5830), .B2(n4837), .C1(n5877), .C2(n5032), .A(n6405), 
        .ZN(n6404) );
  AOI22_X1 U4382 ( .A1(n5879), .A2(n5242), .B1(n5880), .B2(n4967), .ZN(n6405)
         );
  OAI221_X1 U4383 ( .B1(n539), .B2(n5881), .C1(n603), .C2(n5882), .A(n6406), 
        .ZN(n6403) );
  AOI22_X1 U4384 ( .A1(n8110), .A2(n5884), .B1(n8046), .B2(n5885), .ZN(n6406)
         );
  OAI221_X1 U4385 ( .B1(n795), .B2(n5819), .C1(n859), .C2(n5886), .A(n6407), 
        .ZN(n6402) );
  AOI22_X1 U4386 ( .A1(n8238), .A2(n5888), .B1(n8174), .B2(n5889), .ZN(n6407)
         );
  OAI221_X1 U4387 ( .B1(n923), .B2(n5890), .C1(n987), .C2(n5891), .A(n6408), 
        .ZN(n6401) );
  AOI222_X1 U4388 ( .A1(n5893), .A2(n4901), .B1(n5894), .B2(n5160), .C1(n5895), 
        .C2(n5499), .ZN(n6408) );
  OAI22_X1 U4389 ( .A1(n7919), .A2(n5870), .B1(n6409), .B2(n5872), .ZN(n8369)
         );
  NOR4_X1 U4390 ( .A1(n6410), .A2(n6411), .A3(n6412), .A4(n6413), .ZN(n6409)
         );
  OAI221_X1 U4391 ( .B1(n5830), .B2(n4836), .C1(n5877), .C2(n5031), .A(n6414), 
        .ZN(n6413) );
  AOI22_X1 U4392 ( .A1(n5879), .A2(n5241), .B1(n5880), .B2(n4966), .ZN(n6414)
         );
  OAI221_X1 U4393 ( .B1(n540), .B2(n5881), .C1(n604), .C2(n5882), .A(n6415), 
        .ZN(n6412) );
  AOI22_X1 U4394 ( .A1(n8111), .A2(n5884), .B1(n8047), .B2(n5885), .ZN(n6415)
         );
  OAI221_X1 U4395 ( .B1(n796), .B2(n5819), .C1(n860), .C2(n5886), .A(n6416), 
        .ZN(n6411) );
  AOI22_X1 U4396 ( .A1(n8239), .A2(n5888), .B1(n8175), .B2(n5889), .ZN(n6416)
         );
  OAI221_X1 U4397 ( .B1(n924), .B2(n5890), .C1(n988), .C2(n5891), .A(n6417), 
        .ZN(n6410) );
  AOI222_X1 U4398 ( .A1(n5893), .A2(n4900), .B1(n5894), .B2(n5159), .C1(n5895), 
        .C2(n5498), .ZN(n6417) );
  OAI22_X1 U4399 ( .A1(n7920), .A2(n5870), .B1(n6418), .B2(n5872), .ZN(n8370)
         );
  NOR4_X1 U4400 ( .A1(n6419), .A2(n6420), .A3(n6421), .A4(n6422), .ZN(n6418)
         );
  OAI221_X1 U4401 ( .B1(n5830), .B2(n4835), .C1(n5877), .C2(n5030), .A(n6423), 
        .ZN(n6422) );
  AOI22_X1 U4402 ( .A1(n5879), .A2(n5240), .B1(n5880), .B2(n4965), .ZN(n6423)
         );
  OAI221_X1 U4403 ( .B1(n541), .B2(n5881), .C1(n605), .C2(n5882), .A(n6424), 
        .ZN(n6421) );
  AOI22_X1 U4404 ( .A1(n8112), .A2(n5884), .B1(n8048), .B2(n5885), .ZN(n6424)
         );
  OAI221_X1 U4405 ( .B1(n797), .B2(n5819), .C1(n861), .C2(n5886), .A(n6425), 
        .ZN(n6420) );
  AOI22_X1 U4406 ( .A1(n8240), .A2(n5888), .B1(n8176), .B2(n5889), .ZN(n6425)
         );
  OAI221_X1 U4407 ( .B1(n925), .B2(n5890), .C1(n989), .C2(n5891), .A(n6426), 
        .ZN(n6419) );
  AOI222_X1 U4408 ( .A1(n5893), .A2(n4899), .B1(n5894), .B2(n5158), .C1(n5895), 
        .C2(n5497), .ZN(n6426) );
  OAI22_X1 U4409 ( .A1(n7921), .A2(n5870), .B1(n6427), .B2(n5872), .ZN(n8371)
         );
  NOR4_X1 U4410 ( .A1(n6428), .A2(n6429), .A3(n6430), .A4(n6431), .ZN(n6427)
         );
  OAI221_X1 U4411 ( .B1(n5830), .B2(n4834), .C1(n5877), .C2(n5029), .A(n6432), 
        .ZN(n6431) );
  AOI22_X1 U4412 ( .A1(n5879), .A2(n5239), .B1(n5880), .B2(n4964), .ZN(n6432)
         );
  OAI221_X1 U4413 ( .B1(n542), .B2(n5881), .C1(n606), .C2(n5882), .A(n6433), 
        .ZN(n6430) );
  AOI22_X1 U4414 ( .A1(n8113), .A2(n5884), .B1(n8049), .B2(n5885), .ZN(n6433)
         );
  OAI221_X1 U4415 ( .B1(n798), .B2(n5819), .C1(n862), .C2(n5886), .A(n6434), 
        .ZN(n6429) );
  AOI22_X1 U4416 ( .A1(n8241), .A2(n5888), .B1(n8177), .B2(n5889), .ZN(n6434)
         );
  OAI221_X1 U4417 ( .B1(n926), .B2(n5890), .C1(n990), .C2(n5891), .A(n6435), 
        .ZN(n6428) );
  AOI222_X1 U4418 ( .A1(n5893), .A2(n4898), .B1(n5894), .B2(n5157), .C1(n5895), 
        .C2(n5496), .ZN(n6435) );
  OAI22_X1 U4419 ( .A1(n7922), .A2(n5870), .B1(n6436), .B2(n5872), .ZN(n8372)
         );
  NOR4_X1 U4420 ( .A1(n6437), .A2(n6438), .A3(n6439), .A4(n6440), .ZN(n6436)
         );
  OAI221_X1 U4421 ( .B1(n5830), .B2(n4833), .C1(n5877), .C2(n5028), .A(n6441), 
        .ZN(n6440) );
  AOI22_X1 U4422 ( .A1(n5879), .A2(n5238), .B1(n5880), .B2(n4963), .ZN(n6441)
         );
  OAI221_X1 U4423 ( .B1(n543), .B2(n5881), .C1(n607), .C2(n5882), .A(n6442), 
        .ZN(n6439) );
  AOI22_X1 U4424 ( .A1(n8114), .A2(n5884), .B1(n8050), .B2(n5885), .ZN(n6442)
         );
  OAI221_X1 U4425 ( .B1(n799), .B2(n5819), .C1(n863), .C2(n5886), .A(n6443), 
        .ZN(n6438) );
  AOI22_X1 U4426 ( .A1(n8242), .A2(n5888), .B1(n8178), .B2(n5889), .ZN(n6443)
         );
  OAI221_X1 U4427 ( .B1(n927), .B2(n5890), .C1(n991), .C2(n5891), .A(n6444), 
        .ZN(n6437) );
  AOI222_X1 U4428 ( .A1(n5893), .A2(n4897), .B1(n5894), .B2(n5156), .C1(n5895), 
        .C2(n5495), .ZN(n6444) );
  OAI22_X1 U4429 ( .A1(n7923), .A2(n5870), .B1(n6445), .B2(n5872), .ZN(n8373)
         );
  NOR4_X1 U4430 ( .A1(n6446), .A2(n6447), .A3(n6448), .A4(n6449), .ZN(n6445)
         );
  OAI221_X1 U4431 ( .B1(n5830), .B2(n4832), .C1(n5877), .C2(n5027), .A(n6450), 
        .ZN(n6449) );
  AOI22_X1 U4432 ( .A1(n5879), .A2(n5237), .B1(n5880), .B2(n4962), .ZN(n6450)
         );
  OAI221_X1 U4433 ( .B1(n544), .B2(n5881), .C1(n608), .C2(n5882), .A(n6451), 
        .ZN(n6448) );
  AOI22_X1 U4434 ( .A1(n8115), .A2(n5884), .B1(n8051), .B2(n5885), .ZN(n6451)
         );
  OAI221_X1 U4435 ( .B1(n800), .B2(n5819), .C1(n864), .C2(n5886), .A(n6452), 
        .ZN(n6447) );
  AOI22_X1 U4436 ( .A1(n8243), .A2(n5888), .B1(n8179), .B2(n5889), .ZN(n6452)
         );
  OAI221_X1 U4437 ( .B1(n928), .B2(n5890), .C1(n992), .C2(n5891), .A(n6453), 
        .ZN(n6446) );
  AOI222_X1 U4438 ( .A1(n5893), .A2(n4896), .B1(n5894), .B2(n5155), .C1(n5895), 
        .C2(n5494), .ZN(n6453) );
  OAI22_X1 U4439 ( .A1(n7924), .A2(n5870), .B1(n6454), .B2(n5872), .ZN(n8374)
         );
  NOR4_X1 U4440 ( .A1(n6456), .A2(n6457), .A3(n6458), .A4(n6459), .ZN(n6454)
         );
  OAI221_X1 U4441 ( .B1(n5830), .B2(n4831), .C1(n5877), .C2(n5026), .A(n6460), 
        .ZN(n6459) );
  AOI22_X1 U4442 ( .A1(n5879), .A2(n5236), .B1(n5880), .B2(n4961), .ZN(n6460)
         );
  OAI221_X1 U4443 ( .B1(n545), .B2(n5881), .C1(n609), .C2(n5882), .A(n6464), 
        .ZN(n6458) );
  AOI22_X1 U4444 ( .A1(n8116), .A2(n5884), .B1(n8052), .B2(n5885), .ZN(n6464)
         );
  OAI221_X1 U4445 ( .B1(n801), .B2(n5819), .C1(n865), .C2(n5886), .A(n6468), 
        .ZN(n6457) );
  AOI22_X1 U4446 ( .A1(n8244), .A2(n5888), .B1(n8180), .B2(n5889), .ZN(n6468)
         );
  OAI221_X1 U4447 ( .B1(n929), .B2(n5890), .C1(n993), .C2(n5891), .A(n6470), 
        .ZN(n6456) );
  AOI222_X1 U4448 ( .A1(n5893), .A2(n4895), .B1(n5894), .B2(n5154), .C1(n5895), 
        .C2(n5493), .ZN(n6470) );
  INV_X1 U4449 ( .A(n6472), .ZN(n6462) );
  INV_X1 U4450 ( .A(n6473), .ZN(n6465) );
  MUX2_X1 U4451 ( .A(n5831), .B(FILL), .S(n6474), .Z(n8375) );
  AOI21_X1 U4452 ( .B1(n6475), .B2(n6476), .A(n6477), .ZN(n6474) );
  OAI22_X1 U4453 ( .A1(n6478), .A2(n6479), .B1(n1330), .B2(n6480), .ZN(n4830)
         );
  OAI22_X1 U4454 ( .A1(n6481), .A2(n6478), .B1(n1328), .B2(n6480), .ZN(n4829)
         );
  OAI22_X1 U4455 ( .A1(n6482), .A2(n6483), .B1(n6484), .B2(n1250), .ZN(n4828)
         );
  INV_X1 U4456 ( .A(N927), .ZN(n6482) );
  AOI21_X1 U4457 ( .B1(n6484), .B2(n6483), .A(n1261), .ZN(n4827) );
  OAI211_X1 U4458 ( .C1(n1260), .C2(n6484), .A(n6485), .B(n6486), .ZN(n4826)
         );
  NAND3_X1 U4459 ( .A1(n6487), .A2(n6488), .A3(N924), .ZN(n6485) );
  OAI211_X1 U4460 ( .C1(n1259), .C2(n6484), .A(n6489), .B(n6486), .ZN(n4825)
         );
  NAND3_X1 U4461 ( .A1(n6490), .A2(n6491), .A3(n6487), .ZN(n6486) );
  NAND3_X1 U4462 ( .A1(n6487), .A2(n6488), .A3(N925), .ZN(n6489) );
  OAI22_X1 U4463 ( .A1(n6492), .A2(n6483), .B1(n6484), .B2(n1258), .ZN(n4824)
         );
  INV_X1 U4464 ( .A(n6493), .ZN(n6484) );
  OAI211_X1 U4465 ( .C1(CALL), .C2(n6494), .A(n6488), .B(n6487), .ZN(n6483) );
  NOR2_X1 U4466 ( .A1(n6493), .A2(RST), .ZN(n6487) );
  NOR2_X1 U4467 ( .A1(n6477), .A2(n6495), .ZN(n6493) );
  NAND2_X1 U4468 ( .A1(n6455), .A2(n6496), .ZN(n6477) );
  NAND4_X1 U4469 ( .A1(n6497), .A2(RET), .A3(n6498), .A4(n6491), .ZN(n6496) );
  NAND4_X1 U4470 ( .A1(n1250), .A2(n1261), .A3(CALL), .A4(n6499), .ZN(n6488)
         );
  NOR3_X1 U4471 ( .A1(SWP[3]), .A2(n1260), .A3(n1259), .ZN(n6499) );
  INV_X1 U4472 ( .A(N926), .ZN(n6492) );
  MUX2_X1 U4473 ( .A(n6500), .B(SPILL), .S(n6501), .Z(n4823) );
  AOI211_X1 U4474 ( .C1(n6476), .C2(SPILL), .A(RST), .B(n6495), .ZN(n6501) );
  AND4_X1 U4475 ( .A1(n6502), .A2(CALL), .A3(n6503), .A4(n6504), .ZN(n6495) );
  AOI221_X1 U4476 ( .B1(n6505), .B2(SWP[4]), .C1(SWP[1]), .C2(CWP[1]), .A(
        n6506), .ZN(n6504) );
  OAI22_X1 U4477 ( .A1(n1258), .A2(n5862), .B1(n1259), .B2(N890), .ZN(n6506)
         );
  AOI21_X1 U4478 ( .B1(n1318), .B2(n5025), .A(n6507), .ZN(n6503) );
  MUX2_X1 U4479 ( .A(n6490), .B(n6508), .S(n6509), .Z(n6502) );
  INV_X1 U4480 ( .A(n6510), .ZN(n6508) );
  OAI221_X1 U4481 ( .B1(SWP[1]), .B2(CWP[1]), .C1(n5025), .C2(n1318), .A(n6511), .ZN(n6510) );
  AOI222_X1 U4482 ( .A1(n1258), .A2(n5862), .B1(n1259), .B2(N890), .C1(n1250), 
        .C2(n5863), .ZN(n6511) );
  INV_X1 U4483 ( .A(n6494), .ZN(n6490) );
  OAI22_X1 U4484 ( .A1(n6512), .A2(n6478), .B1(n6480), .B2(n5300), .ZN(n4822)
         );
  NAND3_X1 U4485 ( .A1(n6480), .A2(n6455), .A3(n6513), .ZN(n6478) );
  NAND2_X1 U4486 ( .A1(n1327), .A2(n6500), .ZN(n6480) );
  INV_X1 U4487 ( .A(n5870), .ZN(n6500) );
  INV_X1 U4488 ( .A(n6514), .ZN(n6512) );
  OAI221_X1 U4489 ( .B1(n6505), .B2(n6515), .C1(n1303), .C2(n6516), .A(n6517), 
        .ZN(n4821) );
  NAND2_X1 U4490 ( .A1(N916), .A2(n6518), .ZN(n6517) );
  INV_X1 U4491 ( .A(n5863), .ZN(n6505) );
  AOI21_X1 U4492 ( .B1(n6519), .B2(n6516), .A(n1318), .ZN(n4820) );
  NOR2_X1 U4493 ( .A1(n6518), .A2(n6520), .ZN(n6519) );
  INV_X1 U4494 ( .A(n6515), .ZN(n6520) );
  MUX2_X1 U4495 ( .A(n6521), .B(n6522), .S(n1317), .Z(n4819) );
  NAND2_X1 U4496 ( .A1(n6523), .A2(n6515), .ZN(n6522) );
  OAI221_X1 U4497 ( .B1(n6523), .B2(n6524), .C1(N914), .C2(n6515), .A(n6525), 
        .ZN(n4818) );
  AOI22_X1 U4498 ( .A1(N914), .A2(n6526), .B1(n6521), .B2(CWP[2]), .ZN(n6525)
         );
  INV_X1 U4499 ( .A(n6516), .ZN(n6521) );
  OAI221_X1 U4500 ( .B1(n6527), .B2(n6515), .C1(n1315), .C2(n6516), .A(n6528), 
        .ZN(n4817) );
  NAND2_X1 U4501 ( .A1(N915), .A2(n6518), .ZN(n6528) );
  AND2_X1 U4502 ( .A1(n6526), .A2(n6524), .ZN(n6518) );
  NAND3_X1 U4503 ( .A1(n1316), .A2(n1317), .A3(n6529), .ZN(n6524) );
  INV_X1 U4504 ( .A(n6523), .ZN(n6526) );
  NAND3_X1 U4505 ( .A1(n6491), .A2(n6455), .A3(n6516), .ZN(n6523) );
  NAND4_X1 U4506 ( .A1(CALL), .A2(n6516), .A3(n6509), .A4(n6455), .ZN(n6515)
         );
  NAND3_X1 U4507 ( .A1(CWP[2]), .A2(CWP[1]), .A3(n6529), .ZN(n6509) );
  AND3_X1 U4508 ( .A1(n1318), .A2(n1315), .A3(n1303), .ZN(n6529) );
  OAI21_X1 U4509 ( .B1(n6530), .B2(n6507), .A(n6455), .ZN(n6516) );
  NOR2_X1 U4510 ( .A1(CALL), .A2(RET), .ZN(n6530) );
  INV_X1 U4511 ( .A(n5862), .ZN(n6527) );
  MUX2_X1 U4512 ( .A(n6531), .B(n8308), .S(n6532), .Z(n4816) );
  MUX2_X1 U4513 ( .A(n6533), .B(n8307), .S(n6532), .Z(n4815) );
  MUX2_X1 U4514 ( .A(n6534), .B(n8306), .S(n6532), .Z(n4814) );
  MUX2_X1 U4515 ( .A(n6535), .B(n8305), .S(n6532), .Z(n4813) );
  MUX2_X1 U4516 ( .A(n6536), .B(n8304), .S(n6532), .Z(n4812) );
  MUX2_X1 U4517 ( .A(n6537), .B(n8303), .S(n6532), .Z(n4811) );
  MUX2_X1 U4518 ( .A(n6538), .B(n8302), .S(n6532), .Z(n4810) );
  MUX2_X1 U4519 ( .A(n6539), .B(n8301), .S(n6532), .Z(n4809) );
  MUX2_X1 U4520 ( .A(n6540), .B(n8300), .S(n6532), .Z(n4808) );
  MUX2_X1 U4521 ( .A(n6541), .B(n8299), .S(n6532), .Z(n4807) );
  MUX2_X1 U4522 ( .A(n6542), .B(n8298), .S(n6532), .Z(n4806) );
  MUX2_X1 U4523 ( .A(n6543), .B(n8297), .S(n6532), .Z(n4805) );
  MUX2_X1 U4524 ( .A(n6544), .B(n8296), .S(n6532), .Z(n4804) );
  MUX2_X1 U4525 ( .A(n6545), .B(n8295), .S(n6532), .Z(n4803) );
  MUX2_X1 U4526 ( .A(n6546), .B(n8294), .S(n6532), .Z(n4802) );
  MUX2_X1 U4527 ( .A(n6547), .B(n8293), .S(n6532), .Z(n4801) );
  MUX2_X1 U4528 ( .A(n6548), .B(n8292), .S(n6532), .Z(n4800) );
  MUX2_X1 U4529 ( .A(n6549), .B(n8291), .S(n6532), .Z(n4799) );
  MUX2_X1 U4530 ( .A(n6550), .B(n8290), .S(n6532), .Z(n4798) );
  MUX2_X1 U4531 ( .A(n6551), .B(n8289), .S(n6532), .Z(n4797) );
  MUX2_X1 U4532 ( .A(n6552), .B(n8288), .S(n6532), .Z(n4796) );
  MUX2_X1 U4533 ( .A(n6553), .B(n8287), .S(n6532), .Z(n4795) );
  MUX2_X1 U4534 ( .A(n6554), .B(n8286), .S(n6532), .Z(n4794) );
  MUX2_X1 U4535 ( .A(n6555), .B(n8285), .S(n6532), .Z(n4793) );
  MUX2_X1 U4536 ( .A(n6556), .B(n8284), .S(n6532), .Z(n4792) );
  MUX2_X1 U4537 ( .A(n6557), .B(n8283), .S(n6532), .Z(n4791) );
  MUX2_X1 U4538 ( .A(n6558), .B(n8282), .S(n6532), .Z(n4790) );
  MUX2_X1 U4539 ( .A(n6559), .B(n8281), .S(n6532), .Z(n4789) );
  MUX2_X1 U4540 ( .A(n6560), .B(n8280), .S(n6532), .Z(n4788) );
  MUX2_X1 U4541 ( .A(n6561), .B(n8279), .S(n6532), .Z(n4787) );
  MUX2_X1 U4542 ( .A(n6562), .B(n8278), .S(n6532), .Z(n4786) );
  MUX2_X1 U4543 ( .A(n6563), .B(n8277), .S(n6532), .Z(n4785) );
  MUX2_X1 U4544 ( .A(n6564), .B(n8276), .S(n6532), .Z(n4784) );
  MUX2_X1 U4545 ( .A(n6565), .B(n8275), .S(n6532), .Z(n4783) );
  MUX2_X1 U4546 ( .A(n6566), .B(n8274), .S(n6532), .Z(n4782) );
  MUX2_X1 U4547 ( .A(n6567), .B(n8273), .S(n6532), .Z(n4781) );
  MUX2_X1 U4548 ( .A(n6568), .B(n8272), .S(n6532), .Z(n4780) );
  MUX2_X1 U4549 ( .A(n6569), .B(n8271), .S(n6532), .Z(n4779) );
  MUX2_X1 U4550 ( .A(n6570), .B(n8270), .S(n6532), .Z(n4778) );
  MUX2_X1 U4551 ( .A(n6571), .B(n8269), .S(n6532), .Z(n4777) );
  MUX2_X1 U4552 ( .A(n6572), .B(n8268), .S(n6532), .Z(n4776) );
  MUX2_X1 U4553 ( .A(n6573), .B(n8267), .S(n6532), .Z(n4775) );
  MUX2_X1 U4554 ( .A(n6574), .B(n8266), .S(n6532), .Z(n4774) );
  MUX2_X1 U4555 ( .A(n6575), .B(n8265), .S(n6532), .Z(n4773) );
  MUX2_X1 U4556 ( .A(n6576), .B(n8264), .S(n6532), .Z(n4772) );
  MUX2_X1 U4557 ( .A(n6577), .B(n8263), .S(n6532), .Z(n4771) );
  MUX2_X1 U4558 ( .A(n6578), .B(n8262), .S(n6532), .Z(n4770) );
  MUX2_X1 U4559 ( .A(n6579), .B(n8261), .S(n6532), .Z(n4769) );
  MUX2_X1 U4560 ( .A(n6580), .B(n8260), .S(n6532), .Z(n4768) );
  MUX2_X1 U4561 ( .A(n6581), .B(n8259), .S(n6532), .Z(n4767) );
  MUX2_X1 U4562 ( .A(n6582), .B(n8258), .S(n6532), .Z(n4766) );
  MUX2_X1 U4563 ( .A(n6583), .B(n8257), .S(n6532), .Z(n4765) );
  MUX2_X1 U4564 ( .A(n6584), .B(n8256), .S(n6532), .Z(n4764) );
  MUX2_X1 U4565 ( .A(n6585), .B(n8255), .S(n6532), .Z(n4763) );
  MUX2_X1 U4566 ( .A(n6586), .B(n8254), .S(n6532), .Z(n4762) );
  MUX2_X1 U4567 ( .A(n6587), .B(n8253), .S(n6532), .Z(n4761) );
  MUX2_X1 U4568 ( .A(n6588), .B(n8252), .S(n6532), .Z(n4760) );
  MUX2_X1 U4569 ( .A(n6589), .B(n8251), .S(n6532), .Z(n4759) );
  MUX2_X1 U4570 ( .A(n6590), .B(n8250), .S(n6532), .Z(n4758) );
  MUX2_X1 U4571 ( .A(n6591), .B(n8249), .S(n6532), .Z(n4757) );
  MUX2_X1 U4572 ( .A(n6592), .B(n8248), .S(n6532), .Z(n4756) );
  MUX2_X1 U4573 ( .A(n6593), .B(n8247), .S(n6532), .Z(n4755) );
  MUX2_X1 U4574 ( .A(n6594), .B(n8246), .S(n6532), .Z(n4754) );
  MUX2_X1 U4575 ( .A(n6595), .B(n8245), .S(n6532), .Z(n4753) );
  NAND3_X1 U4576 ( .A1(n6598), .A2(n6599), .A3(n6600), .ZN(n6597) );
  NAND4_X1 U4577 ( .A1(n6475), .A2(n5860), .A3(n6461), .A4(n6467), .ZN(n6596)
         );
  MUX2_X1 U4578 ( .A(n5493), .B(n6531), .S(n5844), .Z(n4752) );
  MUX2_X1 U4579 ( .A(n5494), .B(n6533), .S(n5844), .Z(n4751) );
  MUX2_X1 U4580 ( .A(n5495), .B(n6534), .S(n5844), .Z(n4750) );
  MUX2_X1 U4581 ( .A(n5496), .B(n6535), .S(n5844), .Z(n4749) );
  MUX2_X1 U4582 ( .A(n5497), .B(n6536), .S(n5844), .Z(n4748) );
  MUX2_X1 U4583 ( .A(n5498), .B(n6537), .S(n5844), .Z(n4747) );
  MUX2_X1 U4584 ( .A(n5499), .B(n6538), .S(n5844), .Z(n4746) );
  MUX2_X1 U4585 ( .A(n5500), .B(n6539), .S(n5844), .Z(n4745) );
  MUX2_X1 U4586 ( .A(n5501), .B(n6540), .S(n5844), .Z(n4744) );
  MUX2_X1 U4587 ( .A(n5502), .B(n6541), .S(n5844), .Z(n4743) );
  MUX2_X1 U4588 ( .A(n5503), .B(n6542), .S(n5844), .Z(n4742) );
  MUX2_X1 U4589 ( .A(n5504), .B(n6543), .S(n5844), .Z(n4741) );
  MUX2_X1 U4590 ( .A(n5505), .B(n6544), .S(n5844), .Z(n4740) );
  MUX2_X1 U4591 ( .A(n5506), .B(n6545), .S(n5844), .Z(n4739) );
  MUX2_X1 U4592 ( .A(n5507), .B(n6546), .S(n5844), .Z(n4738) );
  MUX2_X1 U4593 ( .A(n5508), .B(n6547), .S(n5844), .Z(n4737) );
  MUX2_X1 U4594 ( .A(n5509), .B(n6548), .S(n5844), .Z(n4736) );
  MUX2_X1 U4595 ( .A(n5510), .B(n6549), .S(n5844), .Z(n4735) );
  MUX2_X1 U4596 ( .A(n5511), .B(n6550), .S(n5844), .Z(n4734) );
  MUX2_X1 U4597 ( .A(n5512), .B(n6551), .S(n5844), .Z(n4733) );
  MUX2_X1 U4598 ( .A(n5513), .B(n6552), .S(n5844), .Z(n4732) );
  MUX2_X1 U4599 ( .A(n5514), .B(n6553), .S(n5844), .Z(n4731) );
  MUX2_X1 U4600 ( .A(n5515), .B(n6554), .S(n5844), .Z(n4730) );
  MUX2_X1 U4601 ( .A(n5516), .B(n6555), .S(n5844), .Z(n4729) );
  MUX2_X1 U4602 ( .A(n5517), .B(n6556), .S(n5844), .Z(n4728) );
  MUX2_X1 U4603 ( .A(n5518), .B(n6557), .S(n5844), .Z(n4727) );
  MUX2_X1 U4604 ( .A(n5519), .B(n6558), .S(n5844), .Z(n4726) );
  MUX2_X1 U4605 ( .A(n5520), .B(n6559), .S(n5844), .Z(n4725) );
  MUX2_X1 U4606 ( .A(n5521), .B(n6560), .S(n5844), .Z(n4724) );
  MUX2_X1 U4607 ( .A(n5522), .B(n6561), .S(n5844), .Z(n4723) );
  MUX2_X1 U4608 ( .A(n5523), .B(n6562), .S(n5844), .Z(n4722) );
  MUX2_X1 U4609 ( .A(n5524), .B(n6563), .S(n5844), .Z(n4721) );
  MUX2_X1 U4610 ( .A(n5525), .B(n6564), .S(n5844), .Z(n4720) );
  MUX2_X1 U4611 ( .A(n5526), .B(n6565), .S(n5844), .Z(n4719) );
  MUX2_X1 U4612 ( .A(n5527), .B(n6566), .S(n5844), .Z(n4718) );
  MUX2_X1 U4613 ( .A(n5528), .B(n6567), .S(n5844), .Z(n4717) );
  MUX2_X1 U4614 ( .A(n5529), .B(n6568), .S(n5844), .Z(n4716) );
  MUX2_X1 U4615 ( .A(n5530), .B(n6569), .S(n5844), .Z(n4715) );
  MUX2_X1 U4616 ( .A(n5531), .B(n6570), .S(n5844), .Z(n4714) );
  MUX2_X1 U4617 ( .A(n5532), .B(n6571), .S(n5844), .Z(n4713) );
  MUX2_X1 U4618 ( .A(n5533), .B(n6572), .S(n5844), .Z(n4712) );
  MUX2_X1 U4619 ( .A(n5534), .B(n6573), .S(n5844), .Z(n4711) );
  MUX2_X1 U4620 ( .A(n5535), .B(n6574), .S(n5844), .Z(n4710) );
  MUX2_X1 U4621 ( .A(n5536), .B(n6575), .S(n5844), .Z(n4709) );
  MUX2_X1 U4622 ( .A(n5537), .B(n6576), .S(n5844), .Z(n4708) );
  MUX2_X1 U4623 ( .A(n5538), .B(n6577), .S(n5844), .Z(n4707) );
  MUX2_X1 U4624 ( .A(n5539), .B(n6578), .S(n5844), .Z(n4706) );
  MUX2_X1 U4625 ( .A(n5540), .B(n6579), .S(n5844), .Z(n4705) );
  MUX2_X1 U4626 ( .A(n5541), .B(n6580), .S(n5844), .Z(n4704) );
  MUX2_X1 U4627 ( .A(n5542), .B(n6581), .S(n5844), .Z(n4703) );
  MUX2_X1 U4628 ( .A(n5543), .B(n6582), .S(n5844), .Z(n4702) );
  MUX2_X1 U4629 ( .A(n5544), .B(n6583), .S(n5844), .Z(n4701) );
  MUX2_X1 U4630 ( .A(n5545), .B(n6584), .S(n5844), .Z(n4700) );
  MUX2_X1 U4631 ( .A(n5546), .B(n6585), .S(n5844), .Z(n4699) );
  MUX2_X1 U4632 ( .A(n5547), .B(n6586), .S(n5844), .Z(n4698) );
  MUX2_X1 U4633 ( .A(n5548), .B(n6587), .S(n5844), .Z(n4697) );
  MUX2_X1 U4634 ( .A(n5549), .B(n6588), .S(n5844), .Z(n4696) );
  MUX2_X1 U4635 ( .A(n5550), .B(n6589), .S(n5844), .Z(n4695) );
  MUX2_X1 U4636 ( .A(n5551), .B(n6590), .S(n5844), .Z(n4694) );
  MUX2_X1 U4637 ( .A(n5552), .B(n6591), .S(n5844), .Z(n4693) );
  MUX2_X1 U4638 ( .A(n5553), .B(n6592), .S(n5844), .Z(n4692) );
  MUX2_X1 U4639 ( .A(n5554), .B(n6593), .S(n5844), .Z(n4691) );
  MUX2_X1 U4640 ( .A(n5555), .B(n6594), .S(n5844), .Z(n4690) );
  MUX2_X1 U4641 ( .A(n5556), .B(n6595), .S(n5844), .Z(n4689) );
  OAI211_X1 U4642 ( .C1(n6473), .C2(n6602), .A(n6603), .B(n6455), .ZN(n6601)
         );
  NAND3_X1 U4643 ( .A1(n6604), .A2(n6605), .A3(n6606), .ZN(n6603) );
  MUX2_X1 U4644 ( .A(n4895), .B(n6531), .S(n5846), .Z(n4688) );
  MUX2_X1 U4645 ( .A(n4896), .B(n6533), .S(n5846), .Z(n4687) );
  MUX2_X1 U4646 ( .A(n4897), .B(n6534), .S(n5846), .Z(n4686) );
  MUX2_X1 U4647 ( .A(n4898), .B(n6535), .S(n5846), .Z(n4685) );
  MUX2_X1 U4648 ( .A(n4899), .B(n6536), .S(n5846), .Z(n4684) );
  MUX2_X1 U4649 ( .A(n4900), .B(n6537), .S(n5846), .Z(n4683) );
  MUX2_X1 U4650 ( .A(n4901), .B(n6538), .S(n5846), .Z(n4682) );
  MUX2_X1 U4651 ( .A(n4902), .B(n6539), .S(n5846), .Z(n4681) );
  MUX2_X1 U4652 ( .A(n4903), .B(n6540), .S(n5846), .Z(n4680) );
  MUX2_X1 U4653 ( .A(n4904), .B(n6541), .S(n5846), .Z(n4679) );
  MUX2_X1 U4654 ( .A(n4905), .B(n6542), .S(n5846), .Z(n4678) );
  MUX2_X1 U4655 ( .A(n4906), .B(n6543), .S(n5846), .Z(n4677) );
  MUX2_X1 U4656 ( .A(n4907), .B(n6544), .S(n5846), .Z(n4676) );
  MUX2_X1 U4657 ( .A(n4908), .B(n6545), .S(n5846), .Z(n4675) );
  MUX2_X1 U4658 ( .A(n4909), .B(n6546), .S(n5846), .Z(n4674) );
  MUX2_X1 U4659 ( .A(n4910), .B(n6547), .S(n5846), .Z(n4673) );
  MUX2_X1 U4660 ( .A(n4911), .B(n6548), .S(n5846), .Z(n4672) );
  MUX2_X1 U4661 ( .A(n4912), .B(n6549), .S(n5846), .Z(n4671) );
  MUX2_X1 U4662 ( .A(n4913), .B(n6550), .S(n5846), .Z(n4670) );
  MUX2_X1 U4663 ( .A(n4914), .B(n6551), .S(n5846), .Z(n4669) );
  MUX2_X1 U4664 ( .A(n4915), .B(n6552), .S(n5846), .Z(n4668) );
  MUX2_X1 U4665 ( .A(n4916), .B(n6553), .S(n5846), .Z(n4667) );
  MUX2_X1 U4666 ( .A(n4917), .B(n6554), .S(n5846), .Z(n4666) );
  MUX2_X1 U4667 ( .A(n4918), .B(n6555), .S(n5846), .Z(n4665) );
  MUX2_X1 U4668 ( .A(n4919), .B(n6556), .S(n5846), .Z(n4664) );
  MUX2_X1 U4669 ( .A(n4920), .B(n6557), .S(n5846), .Z(n4663) );
  MUX2_X1 U4670 ( .A(n4921), .B(n6558), .S(n5846), .Z(n4662) );
  MUX2_X1 U4671 ( .A(n4922), .B(n6559), .S(n5846), .Z(n4661) );
  MUX2_X1 U4672 ( .A(n4923), .B(n6560), .S(n5846), .Z(n4660) );
  MUX2_X1 U4673 ( .A(n4924), .B(n6561), .S(n5846), .Z(n4659) );
  MUX2_X1 U4674 ( .A(n4925), .B(n6562), .S(n5846), .Z(n4658) );
  MUX2_X1 U4675 ( .A(n4926), .B(n6563), .S(n5846), .Z(n4657) );
  MUX2_X1 U4676 ( .A(n4927), .B(n6564), .S(n5846), .Z(n4656) );
  MUX2_X1 U4677 ( .A(n4928), .B(n6565), .S(n5846), .Z(n4655) );
  MUX2_X1 U4678 ( .A(n4929), .B(n6566), .S(n5846), .Z(n4654) );
  MUX2_X1 U4679 ( .A(n4930), .B(n6567), .S(n5846), .Z(n4653) );
  MUX2_X1 U4680 ( .A(n4931), .B(n6568), .S(n5846), .Z(n4652) );
  MUX2_X1 U4681 ( .A(n4932), .B(n6569), .S(n5846), .Z(n4651) );
  MUX2_X1 U4682 ( .A(n4933), .B(n6570), .S(n5846), .Z(n4650) );
  MUX2_X1 U4683 ( .A(n4934), .B(n6571), .S(n5846), .Z(n4649) );
  MUX2_X1 U4684 ( .A(n4935), .B(n6572), .S(n5846), .Z(n4648) );
  MUX2_X1 U4685 ( .A(n4936), .B(n6573), .S(n5846), .Z(n4647) );
  MUX2_X1 U4686 ( .A(n4937), .B(n6574), .S(n5846), .Z(n4646) );
  MUX2_X1 U4687 ( .A(n4938), .B(n6575), .S(n5846), .Z(n4645) );
  MUX2_X1 U4688 ( .A(n4939), .B(n6576), .S(n5846), .Z(n4644) );
  MUX2_X1 U4689 ( .A(n4940), .B(n6577), .S(n5846), .Z(n4643) );
  MUX2_X1 U4690 ( .A(n4941), .B(n6578), .S(n5846), .Z(n4642) );
  MUX2_X1 U4691 ( .A(n4942), .B(n6579), .S(n5846), .Z(n4641) );
  MUX2_X1 U4692 ( .A(n4943), .B(n6580), .S(n5846), .Z(n4640) );
  MUX2_X1 U4693 ( .A(n4944), .B(n6581), .S(n5846), .Z(n4639) );
  MUX2_X1 U4694 ( .A(n4945), .B(n6582), .S(n5846), .Z(n4638) );
  MUX2_X1 U4695 ( .A(n4946), .B(n6583), .S(n5846), .Z(n4637) );
  MUX2_X1 U4696 ( .A(n4947), .B(n6584), .S(n5846), .Z(n4636) );
  MUX2_X1 U4697 ( .A(n4948), .B(n6585), .S(n5846), .Z(n4635) );
  MUX2_X1 U4698 ( .A(n4949), .B(n6586), .S(n5846), .Z(n4634) );
  MUX2_X1 U4699 ( .A(n4950), .B(n6587), .S(n5846), .Z(n4633) );
  MUX2_X1 U4700 ( .A(n4951), .B(n6588), .S(n5846), .Z(n4632) );
  MUX2_X1 U4701 ( .A(n4952), .B(n6589), .S(n5846), .Z(n4631) );
  MUX2_X1 U4702 ( .A(n4953), .B(n6590), .S(n5846), .Z(n4630) );
  MUX2_X1 U4703 ( .A(n4954), .B(n6591), .S(n5846), .Z(n4629) );
  MUX2_X1 U4704 ( .A(n4955), .B(n6592), .S(n5846), .Z(n4628) );
  MUX2_X1 U4705 ( .A(n4956), .B(n6593), .S(n5846), .Z(n4627) );
  MUX2_X1 U4706 ( .A(n4957), .B(n6594), .S(n5846), .Z(n4626) );
  MUX2_X1 U4707 ( .A(n4958), .B(n6595), .S(n5846), .Z(n4625) );
  OAI211_X1 U4708 ( .C1(n6472), .C2(n6602), .A(n6608), .B(n6455), .ZN(n6607)
         );
  NAND3_X1 U4709 ( .A1(n6606), .A2(n6609), .A3(n6610), .ZN(n6608) );
  MUX2_X1 U4710 ( .A(n6531), .B(n5154), .S(n6611), .Z(n4624) );
  MUX2_X1 U4711 ( .A(n6533), .B(n5155), .S(n6611), .Z(n4623) );
  MUX2_X1 U4712 ( .A(n6534), .B(n5156), .S(n6611), .Z(n4622) );
  MUX2_X1 U4713 ( .A(n6535), .B(n5157), .S(n6611), .Z(n4621) );
  MUX2_X1 U4714 ( .A(n6536), .B(n5158), .S(n6611), .Z(n4620) );
  MUX2_X1 U4715 ( .A(n6537), .B(n5159), .S(n6611), .Z(n4619) );
  MUX2_X1 U4716 ( .A(n6538), .B(n5160), .S(n6611), .Z(n4618) );
  MUX2_X1 U4717 ( .A(n6539), .B(n5161), .S(n6611), .Z(n4617) );
  MUX2_X1 U4718 ( .A(n6540), .B(n5162), .S(n6611), .Z(n4616) );
  MUX2_X1 U4719 ( .A(n6541), .B(n5163), .S(n6611), .Z(n4615) );
  MUX2_X1 U4720 ( .A(n6542), .B(n5164), .S(n6611), .Z(n4614) );
  MUX2_X1 U4721 ( .A(n6543), .B(n5165), .S(n6611), .Z(n4613) );
  MUX2_X1 U4722 ( .A(n6544), .B(n5166), .S(n6611), .Z(n4612) );
  MUX2_X1 U4723 ( .A(n6545), .B(n5167), .S(n6611), .Z(n4611) );
  MUX2_X1 U4724 ( .A(n6546), .B(n5168), .S(n6611), .Z(n4610) );
  MUX2_X1 U4725 ( .A(n6547), .B(n5169), .S(n6611), .Z(n4609) );
  MUX2_X1 U4726 ( .A(n6548), .B(n5170), .S(n6611), .Z(n4608) );
  MUX2_X1 U4727 ( .A(n6549), .B(n5171), .S(n6611), .Z(n4607) );
  MUX2_X1 U4728 ( .A(n6550), .B(n5172), .S(n6611), .Z(n4606) );
  MUX2_X1 U4729 ( .A(n6551), .B(n5173), .S(n6611), .Z(n4605) );
  MUX2_X1 U4730 ( .A(n6552), .B(n5174), .S(n6611), .Z(n4604) );
  MUX2_X1 U4731 ( .A(n6553), .B(n5175), .S(n6611), .Z(n4603) );
  MUX2_X1 U4732 ( .A(n6554), .B(n5176), .S(n6611), .Z(n4602) );
  MUX2_X1 U4733 ( .A(n6555), .B(n5177), .S(n6611), .Z(n4601) );
  MUX2_X1 U4734 ( .A(n6556), .B(n5178), .S(n6611), .Z(n4600) );
  MUX2_X1 U4735 ( .A(n6557), .B(n5179), .S(n6611), .Z(n4599) );
  MUX2_X1 U4736 ( .A(n6558), .B(n5180), .S(n6611), .Z(n4598) );
  MUX2_X1 U4737 ( .A(n6559), .B(n5181), .S(n6611), .Z(n4597) );
  MUX2_X1 U4738 ( .A(n6560), .B(n5182), .S(n6611), .Z(n4596) );
  MUX2_X1 U4739 ( .A(n6561), .B(n5183), .S(n6611), .Z(n4595) );
  MUX2_X1 U4740 ( .A(n6562), .B(n5184), .S(n6611), .Z(n4594) );
  MUX2_X1 U4741 ( .A(n6563), .B(n5185), .S(n6611), .Z(n4593) );
  MUX2_X1 U4742 ( .A(n6564), .B(n5186), .S(n6611), .Z(n4592) );
  MUX2_X1 U4743 ( .A(n6565), .B(n5187), .S(n6611), .Z(n4591) );
  MUX2_X1 U4744 ( .A(n6566), .B(n5188), .S(n6611), .Z(n4590) );
  MUX2_X1 U4745 ( .A(n6567), .B(n5189), .S(n6611), .Z(n4589) );
  MUX2_X1 U4746 ( .A(n6568), .B(n5190), .S(n6611), .Z(n4588) );
  MUX2_X1 U4747 ( .A(n6569), .B(n5191), .S(n6611), .Z(n4587) );
  MUX2_X1 U4748 ( .A(n6570), .B(n5192), .S(n6611), .Z(n4586) );
  MUX2_X1 U4749 ( .A(n6571), .B(n5193), .S(n6611), .Z(n4585) );
  MUX2_X1 U4750 ( .A(n6572), .B(n5194), .S(n6611), .Z(n4584) );
  MUX2_X1 U4751 ( .A(n6573), .B(n5195), .S(n6611), .Z(n4583) );
  MUX2_X1 U4752 ( .A(n6574), .B(n5196), .S(n6611), .Z(n4582) );
  MUX2_X1 U4753 ( .A(n6575), .B(n5197), .S(n6611), .Z(n4581) );
  MUX2_X1 U4754 ( .A(n6576), .B(n5198), .S(n6611), .Z(n4580) );
  MUX2_X1 U4755 ( .A(n6577), .B(n5199), .S(n6611), .Z(n4579) );
  MUX2_X1 U4756 ( .A(n6578), .B(n5200), .S(n6611), .Z(n4578) );
  MUX2_X1 U4757 ( .A(n6579), .B(n5201), .S(n6611), .Z(n4577) );
  MUX2_X1 U4758 ( .A(n6580), .B(n5202), .S(n6611), .Z(n4576) );
  MUX2_X1 U4759 ( .A(n6581), .B(n5203), .S(n6611), .Z(n4575) );
  MUX2_X1 U4760 ( .A(n6582), .B(n5204), .S(n6611), .Z(n4574) );
  MUX2_X1 U4761 ( .A(n6583), .B(n5205), .S(n6611), .Z(n4573) );
  MUX2_X1 U4762 ( .A(n6584), .B(n5206), .S(n6611), .Z(n4572) );
  MUX2_X1 U4763 ( .A(n6585), .B(n5207), .S(n6611), .Z(n4571) );
  MUX2_X1 U4764 ( .A(n6586), .B(n5208), .S(n6611), .Z(n4570) );
  MUX2_X1 U4765 ( .A(n6587), .B(n5209), .S(n6611), .Z(n4569) );
  MUX2_X1 U4766 ( .A(n6588), .B(n5210), .S(n6611), .Z(n4568) );
  MUX2_X1 U4767 ( .A(n6589), .B(n5211), .S(n6611), .Z(n4567) );
  MUX2_X1 U4768 ( .A(n6590), .B(n5212), .S(n6611), .Z(n4566) );
  MUX2_X1 U4769 ( .A(n6591), .B(n5213), .S(n6611), .Z(n4565) );
  MUX2_X1 U4770 ( .A(n6592), .B(n5214), .S(n6611), .Z(n4564) );
  MUX2_X1 U4771 ( .A(n6593), .B(n5215), .S(n6611), .Z(n4563) );
  MUX2_X1 U4772 ( .A(n6594), .B(n5216), .S(n6611), .Z(n4562) );
  MUX2_X1 U4773 ( .A(n6595), .B(n5217), .S(n6611), .Z(n4561) );
  MUX2_X1 U4774 ( .A(n6531), .B(n5687), .S(n6614), .Z(n4560) );
  MUX2_X1 U4775 ( .A(n6533), .B(n5688), .S(n6614), .Z(n4559) );
  MUX2_X1 U4776 ( .A(n6534), .B(n5689), .S(n6614), .Z(n4558) );
  MUX2_X1 U4777 ( .A(n6535), .B(n5690), .S(n6614), .Z(n4557) );
  MUX2_X1 U4778 ( .A(n6536), .B(n5691), .S(n6614), .Z(n4556) );
  MUX2_X1 U4779 ( .A(n6537), .B(n5692), .S(n6614), .Z(n4555) );
  MUX2_X1 U4780 ( .A(n6538), .B(n5693), .S(n6614), .Z(n4554) );
  MUX2_X1 U4781 ( .A(n6539), .B(n5694), .S(n6614), .Z(n4553) );
  MUX2_X1 U4782 ( .A(n6540), .B(n5695), .S(n6614), .Z(n4552) );
  MUX2_X1 U4783 ( .A(n6541), .B(n5696), .S(n6614), .Z(n4551) );
  MUX2_X1 U4784 ( .A(n6542), .B(n5697), .S(n6614), .Z(n4550) );
  MUX2_X1 U4785 ( .A(n6543), .B(n5698), .S(n6614), .Z(n4549) );
  MUX2_X1 U4786 ( .A(n6544), .B(n5699), .S(n6614), .Z(n4548) );
  MUX2_X1 U4787 ( .A(n6545), .B(n5700), .S(n6614), .Z(n4547) );
  MUX2_X1 U4788 ( .A(n6546), .B(n5701), .S(n6614), .Z(n4546) );
  MUX2_X1 U4789 ( .A(n6547), .B(n5702), .S(n6614), .Z(n4545) );
  MUX2_X1 U4790 ( .A(n6548), .B(n5703), .S(n6614), .Z(n4544) );
  MUX2_X1 U4791 ( .A(n6549), .B(n5704), .S(n6614), .Z(n4543) );
  MUX2_X1 U4792 ( .A(n6550), .B(n5705), .S(n6614), .Z(n4542) );
  MUX2_X1 U4793 ( .A(n6551), .B(n5706), .S(n6614), .Z(n4541) );
  MUX2_X1 U4794 ( .A(n6552), .B(n5707), .S(n6614), .Z(n4540) );
  MUX2_X1 U4795 ( .A(n6553), .B(n5708), .S(n6614), .Z(n4539) );
  MUX2_X1 U4796 ( .A(n6554), .B(n5709), .S(n6614), .Z(n4538) );
  MUX2_X1 U4797 ( .A(n6555), .B(n5710), .S(n6614), .Z(n4537) );
  MUX2_X1 U4798 ( .A(n6556), .B(n5711), .S(n6614), .Z(n4536) );
  MUX2_X1 U4799 ( .A(n6557), .B(n5712), .S(n6614), .Z(n4535) );
  MUX2_X1 U4800 ( .A(n6558), .B(n5713), .S(n6614), .Z(n4534) );
  MUX2_X1 U4801 ( .A(n6559), .B(n5714), .S(n6614), .Z(n4533) );
  MUX2_X1 U4802 ( .A(n6560), .B(n5715), .S(n6614), .Z(n4532) );
  MUX2_X1 U4803 ( .A(n6561), .B(n5716), .S(n6614), .Z(n4531) );
  MUX2_X1 U4804 ( .A(n6562), .B(n5717), .S(n6614), .Z(n4530) );
  MUX2_X1 U4805 ( .A(n6563), .B(n5718), .S(n6614), .Z(n4529) );
  MUX2_X1 U4806 ( .A(n6564), .B(n5719), .S(n6614), .Z(n4528) );
  MUX2_X1 U4807 ( .A(n6565), .B(n5720), .S(n6614), .Z(n4527) );
  MUX2_X1 U4808 ( .A(n6566), .B(n5721), .S(n6614), .Z(n4526) );
  MUX2_X1 U4809 ( .A(n6567), .B(n5722), .S(n6614), .Z(n4525) );
  MUX2_X1 U4810 ( .A(n6568), .B(n5723), .S(n6614), .Z(n4524) );
  MUX2_X1 U4811 ( .A(n6569), .B(n5724), .S(n6614), .Z(n4523) );
  MUX2_X1 U4812 ( .A(n6570), .B(n5725), .S(n6614), .Z(n4522) );
  MUX2_X1 U4813 ( .A(n6571), .B(n5726), .S(n6614), .Z(n4521) );
  MUX2_X1 U4814 ( .A(n6572), .B(n5727), .S(n6614), .Z(n4520) );
  MUX2_X1 U4815 ( .A(n6573), .B(n5728), .S(n6614), .Z(n4519) );
  MUX2_X1 U4816 ( .A(n6574), .B(n5729), .S(n6614), .Z(n4518) );
  MUX2_X1 U4817 ( .A(n6575), .B(n5730), .S(n6614), .Z(n4517) );
  MUX2_X1 U4818 ( .A(n6576), .B(n5731), .S(n6614), .Z(n4516) );
  MUX2_X1 U4819 ( .A(n6577), .B(n5732), .S(n6614), .Z(n4515) );
  MUX2_X1 U4820 ( .A(n6578), .B(n5733), .S(n6614), .Z(n4514) );
  MUX2_X1 U4821 ( .A(n6579), .B(n5734), .S(n6614), .Z(n4513) );
  MUX2_X1 U4822 ( .A(n6580), .B(n5735), .S(n6614), .Z(n4512) );
  MUX2_X1 U4823 ( .A(n6581), .B(n5736), .S(n6614), .Z(n4511) );
  MUX2_X1 U4824 ( .A(n6582), .B(n5737), .S(n6614), .Z(n4510) );
  MUX2_X1 U4825 ( .A(n6583), .B(n5738), .S(n6614), .Z(n4509) );
  MUX2_X1 U4826 ( .A(n6584), .B(n5739), .S(n6614), .Z(n4508) );
  MUX2_X1 U4827 ( .A(n6585), .B(n5740), .S(n6614), .Z(n4507) );
  MUX2_X1 U4828 ( .A(n6586), .B(n5741), .S(n6614), .Z(n4506) );
  MUX2_X1 U4829 ( .A(n6587), .B(n5742), .S(n6614), .Z(n4505) );
  MUX2_X1 U4830 ( .A(n6588), .B(n5743), .S(n6614), .Z(n4504) );
  MUX2_X1 U4831 ( .A(n6589), .B(n5744), .S(n6614), .Z(n4503) );
  MUX2_X1 U4832 ( .A(n6590), .B(n5745), .S(n6614), .Z(n4502) );
  MUX2_X1 U4833 ( .A(n6591), .B(n5746), .S(n6614), .Z(n4501) );
  MUX2_X1 U4834 ( .A(n6592), .B(n5747), .S(n6614), .Z(n4500) );
  MUX2_X1 U4835 ( .A(n6593), .B(n5748), .S(n6614), .Z(n4499) );
  MUX2_X1 U4836 ( .A(n6594), .B(n5749), .S(n6614), .Z(n4498) );
  MUX2_X1 U4837 ( .A(n6595), .B(n5750), .S(n6614), .Z(n4497) );
  AND3_X1 U4838 ( .A1(n6609), .A2(n6616), .A3(n6612), .ZN(n6615) );
  INV_X1 U4839 ( .A(n6602), .ZN(n6613) );
  NAND2_X1 U4840 ( .A1(n6617), .A2(n6471), .ZN(n6602) );
  NOR2_X1 U4841 ( .A1(n6618), .A2(n6619), .ZN(n6471) );
  MUX2_X1 U4842 ( .A(n5090), .B(n6531), .S(n5848), .Z(n4496) );
  MUX2_X1 U4843 ( .A(n5091), .B(n6533), .S(n5848), .Z(n4495) );
  MUX2_X1 U4844 ( .A(n5092), .B(n6534), .S(n5848), .Z(n4494) );
  MUX2_X1 U4845 ( .A(n5093), .B(n6535), .S(n5848), .Z(n4493) );
  MUX2_X1 U4846 ( .A(n5094), .B(n6536), .S(n5848), .Z(n4492) );
  MUX2_X1 U4847 ( .A(n5095), .B(n6537), .S(n5848), .Z(n4491) );
  MUX2_X1 U4848 ( .A(n5096), .B(n6538), .S(n5848), .Z(n4490) );
  MUX2_X1 U4849 ( .A(n5097), .B(n6539), .S(n5848), .Z(n4489) );
  MUX2_X1 U4850 ( .A(n5098), .B(n6540), .S(n5848), .Z(n4488) );
  MUX2_X1 U4851 ( .A(n5099), .B(n6541), .S(n5848), .Z(n4487) );
  MUX2_X1 U4852 ( .A(n5100), .B(n6542), .S(n5848), .Z(n4486) );
  MUX2_X1 U4853 ( .A(n5101), .B(n6543), .S(n5848), .Z(n4485) );
  MUX2_X1 U4854 ( .A(n5102), .B(n6544), .S(n5848), .Z(n4484) );
  MUX2_X1 U4855 ( .A(n5103), .B(n6545), .S(n5848), .Z(n4483) );
  MUX2_X1 U4856 ( .A(n5104), .B(n6546), .S(n5848), .Z(n4482) );
  MUX2_X1 U4857 ( .A(n5105), .B(n6547), .S(n5848), .Z(n4481) );
  MUX2_X1 U4858 ( .A(n5106), .B(n6548), .S(n5848), .Z(n4480) );
  MUX2_X1 U4859 ( .A(n5107), .B(n6549), .S(n5848), .Z(n4479) );
  MUX2_X1 U4860 ( .A(n5108), .B(n6550), .S(n5848), .Z(n4478) );
  MUX2_X1 U4861 ( .A(n5109), .B(n6551), .S(n5848), .Z(n4477) );
  MUX2_X1 U4862 ( .A(n5110), .B(n6552), .S(n5848), .Z(n4476) );
  MUX2_X1 U4863 ( .A(n5111), .B(n6553), .S(n5848), .Z(n4475) );
  MUX2_X1 U4864 ( .A(n5112), .B(n6554), .S(n5848), .Z(n4474) );
  MUX2_X1 U4865 ( .A(n5113), .B(n6555), .S(n5848), .Z(n4473) );
  MUX2_X1 U4866 ( .A(n5114), .B(n6556), .S(n5848), .Z(n4472) );
  MUX2_X1 U4867 ( .A(n5115), .B(n6557), .S(n5848), .Z(n4471) );
  MUX2_X1 U4868 ( .A(n5116), .B(n6558), .S(n5848), .Z(n4470) );
  MUX2_X1 U4869 ( .A(n5117), .B(n6559), .S(n5848), .Z(n4469) );
  MUX2_X1 U4870 ( .A(n5118), .B(n6560), .S(n5848), .Z(n4468) );
  MUX2_X1 U4871 ( .A(n5119), .B(n6561), .S(n5848), .Z(n4467) );
  MUX2_X1 U4872 ( .A(n5120), .B(n6562), .S(n5848), .Z(n4466) );
  MUX2_X1 U4873 ( .A(n5121), .B(n6563), .S(n5848), .Z(n4465) );
  MUX2_X1 U4874 ( .A(n5122), .B(n6564), .S(n5848), .Z(n4464) );
  MUX2_X1 U4875 ( .A(n5123), .B(n6565), .S(n5848), .Z(n4463) );
  MUX2_X1 U4876 ( .A(n5124), .B(n6566), .S(n5848), .Z(n4462) );
  MUX2_X1 U4877 ( .A(n5125), .B(n6567), .S(n5848), .Z(n4461) );
  MUX2_X1 U4878 ( .A(n5126), .B(n6568), .S(n5848), .Z(n4460) );
  MUX2_X1 U4879 ( .A(n5127), .B(n6569), .S(n5848), .Z(n4459) );
  MUX2_X1 U4880 ( .A(n5128), .B(n6570), .S(n5848), .Z(n4458) );
  MUX2_X1 U4881 ( .A(n5129), .B(n6571), .S(n5848), .Z(n4457) );
  MUX2_X1 U4882 ( .A(n5130), .B(n6572), .S(n5848), .Z(n4456) );
  MUX2_X1 U4883 ( .A(n5131), .B(n6573), .S(n5848), .Z(n4455) );
  MUX2_X1 U4884 ( .A(n5132), .B(n6574), .S(n5848), .Z(n4454) );
  MUX2_X1 U4885 ( .A(n5133), .B(n6575), .S(n5848), .Z(n4453) );
  MUX2_X1 U4886 ( .A(n5134), .B(n6576), .S(n5848), .Z(n4452) );
  MUX2_X1 U4887 ( .A(n5135), .B(n6577), .S(n5848), .Z(n4451) );
  MUX2_X1 U4888 ( .A(n5136), .B(n6578), .S(n5848), .Z(n4450) );
  MUX2_X1 U4889 ( .A(n5137), .B(n6579), .S(n5848), .Z(n4449) );
  MUX2_X1 U4890 ( .A(n5138), .B(n6580), .S(n5848), .Z(n4448) );
  MUX2_X1 U4891 ( .A(n5139), .B(n6581), .S(n5848), .Z(n4447) );
  MUX2_X1 U4892 ( .A(n5140), .B(n6582), .S(n5848), .Z(n4446) );
  MUX2_X1 U4893 ( .A(n5141), .B(n6583), .S(n5848), .Z(n4445) );
  MUX2_X1 U4894 ( .A(n5142), .B(n6584), .S(n5848), .Z(n4444) );
  MUX2_X1 U4895 ( .A(n5143), .B(n6585), .S(n5848), .Z(n4443) );
  MUX2_X1 U4896 ( .A(n5144), .B(n6586), .S(n5848), .Z(n4442) );
  MUX2_X1 U4897 ( .A(n5145), .B(n6587), .S(n5848), .Z(n4441) );
  MUX2_X1 U4898 ( .A(n5146), .B(n6588), .S(n5848), .Z(n4440) );
  MUX2_X1 U4899 ( .A(n5147), .B(n6589), .S(n5848), .Z(n4439) );
  MUX2_X1 U4900 ( .A(n5148), .B(n6590), .S(n5848), .Z(n4438) );
  MUX2_X1 U4901 ( .A(n5149), .B(n6591), .S(n5848), .Z(n4437) );
  MUX2_X1 U4902 ( .A(n5150), .B(n6592), .S(n5848), .Z(n4436) );
  MUX2_X1 U4903 ( .A(n5151), .B(n6593), .S(n5848), .Z(n4435) );
  MUX2_X1 U4904 ( .A(n5152), .B(n6594), .S(n5848), .Z(n4434) );
  MUX2_X1 U4905 ( .A(n5153), .B(n6595), .S(n5848), .Z(n4433) );
  OAI211_X1 U4906 ( .C1(n6473), .C2(n6621), .A(n6622), .B(n6455), .ZN(n6620)
         );
  NAND3_X1 U4907 ( .A1(n6604), .A2(n6623), .A3(n6605), .ZN(n6622) );
  MUX2_X1 U4908 ( .A(n5301), .B(n6531), .S(n5850), .Z(n4432) );
  MUX2_X1 U4909 ( .A(n5302), .B(n6533), .S(n5850), .Z(n4431) );
  MUX2_X1 U4910 ( .A(n5303), .B(n6534), .S(n5850), .Z(n4430) );
  MUX2_X1 U4911 ( .A(n5304), .B(n6535), .S(n5850), .Z(n4429) );
  MUX2_X1 U4912 ( .A(n5305), .B(n6536), .S(n5850), .Z(n4428) );
  MUX2_X1 U4913 ( .A(n5306), .B(n6537), .S(n5850), .Z(n4427) );
  MUX2_X1 U4914 ( .A(n5307), .B(n6538), .S(n5850), .Z(n4426) );
  MUX2_X1 U4915 ( .A(n5308), .B(n6539), .S(n5850), .Z(n4425) );
  MUX2_X1 U4916 ( .A(n5309), .B(n6540), .S(n5850), .Z(n4424) );
  MUX2_X1 U4917 ( .A(n5310), .B(n6541), .S(n5850), .Z(n4423) );
  MUX2_X1 U4918 ( .A(n5311), .B(n6542), .S(n5850), .Z(n4422) );
  MUX2_X1 U4919 ( .A(n5312), .B(n6543), .S(n5850), .Z(n4421) );
  MUX2_X1 U4920 ( .A(n5313), .B(n6544), .S(n5850), .Z(n4420) );
  MUX2_X1 U4921 ( .A(n5314), .B(n6545), .S(n5850), .Z(n4419) );
  MUX2_X1 U4922 ( .A(n5315), .B(n6546), .S(n5850), .Z(n4418) );
  MUX2_X1 U4923 ( .A(n5316), .B(n6547), .S(n5850), .Z(n4417) );
  MUX2_X1 U4924 ( .A(n5317), .B(n6548), .S(n5850), .Z(n4416) );
  MUX2_X1 U4925 ( .A(n5318), .B(n6549), .S(n5850), .Z(n4415) );
  MUX2_X1 U4926 ( .A(n5319), .B(n6550), .S(n5850), .Z(n4414) );
  MUX2_X1 U4927 ( .A(n5320), .B(n6551), .S(n5850), .Z(n4413) );
  MUX2_X1 U4928 ( .A(n5321), .B(n6552), .S(n5850), .Z(n4412) );
  MUX2_X1 U4929 ( .A(n5322), .B(n6553), .S(n5850), .Z(n4411) );
  MUX2_X1 U4930 ( .A(n5323), .B(n6554), .S(n5850), .Z(n4410) );
  MUX2_X1 U4931 ( .A(n5324), .B(n6555), .S(n5850), .Z(n4409) );
  MUX2_X1 U4932 ( .A(n5325), .B(n6556), .S(n5850), .Z(n4408) );
  MUX2_X1 U4933 ( .A(n5326), .B(n6557), .S(n5850), .Z(n4407) );
  MUX2_X1 U4934 ( .A(n5327), .B(n6558), .S(n5850), .Z(n4406) );
  MUX2_X1 U4935 ( .A(n5328), .B(n6559), .S(n5850), .Z(n4405) );
  MUX2_X1 U4936 ( .A(n5329), .B(n6560), .S(n5850), .Z(n4404) );
  MUX2_X1 U4937 ( .A(n5330), .B(n6561), .S(n5850), .Z(n4403) );
  MUX2_X1 U4938 ( .A(n5331), .B(n6562), .S(n5850), .Z(n4402) );
  MUX2_X1 U4939 ( .A(n5332), .B(n6563), .S(n5850), .Z(n4401) );
  MUX2_X1 U4940 ( .A(n5333), .B(n6564), .S(n5850), .Z(n4400) );
  MUX2_X1 U4941 ( .A(n5334), .B(n6565), .S(n5850), .Z(n4399) );
  MUX2_X1 U4942 ( .A(n5335), .B(n6566), .S(n5850), .Z(n4398) );
  MUX2_X1 U4943 ( .A(n5336), .B(n6567), .S(n5850), .Z(n4397) );
  MUX2_X1 U4944 ( .A(n5337), .B(n6568), .S(n5850), .Z(n4396) );
  MUX2_X1 U4945 ( .A(n5338), .B(n6569), .S(n5850), .Z(n4395) );
  MUX2_X1 U4946 ( .A(n5339), .B(n6570), .S(n5850), .Z(n4394) );
  MUX2_X1 U4947 ( .A(n5340), .B(n6571), .S(n5850), .Z(n4393) );
  MUX2_X1 U4948 ( .A(n5341), .B(n6572), .S(n5850), .Z(n4392) );
  MUX2_X1 U4949 ( .A(n5342), .B(n6573), .S(n5850), .Z(n4391) );
  MUX2_X1 U4950 ( .A(n5343), .B(n6574), .S(n5850), .Z(n4390) );
  MUX2_X1 U4951 ( .A(n5344), .B(n6575), .S(n5850), .Z(n4389) );
  MUX2_X1 U4952 ( .A(n5345), .B(n6576), .S(n5850), .Z(n4388) );
  MUX2_X1 U4953 ( .A(n5346), .B(n6577), .S(n5850), .Z(n4387) );
  MUX2_X1 U4954 ( .A(n5347), .B(n6578), .S(n5850), .Z(n4386) );
  MUX2_X1 U4955 ( .A(n5348), .B(n6579), .S(n5850), .Z(n4385) );
  MUX2_X1 U4956 ( .A(n5349), .B(n6580), .S(n5850), .Z(n4384) );
  MUX2_X1 U4957 ( .A(n5350), .B(n6581), .S(n5850), .Z(n4383) );
  MUX2_X1 U4958 ( .A(n5351), .B(n6582), .S(n5850), .Z(n4382) );
  MUX2_X1 U4959 ( .A(n5352), .B(n6583), .S(n5850), .Z(n4381) );
  MUX2_X1 U4960 ( .A(n5353), .B(n6584), .S(n5850), .Z(n4380) );
  MUX2_X1 U4961 ( .A(n5354), .B(n6585), .S(n5850), .Z(n4379) );
  MUX2_X1 U4962 ( .A(n5355), .B(n6586), .S(n5850), .Z(n4378) );
  MUX2_X1 U4963 ( .A(n5356), .B(n6587), .S(n5850), .Z(n4377) );
  MUX2_X1 U4964 ( .A(n5357), .B(n6588), .S(n5850), .Z(n4376) );
  MUX2_X1 U4965 ( .A(n5358), .B(n6589), .S(n5850), .Z(n4375) );
  MUX2_X1 U4966 ( .A(n5359), .B(n6590), .S(n5850), .Z(n4374) );
  MUX2_X1 U4967 ( .A(n5360), .B(n6591), .S(n5850), .Z(n4373) );
  MUX2_X1 U4968 ( .A(n5361), .B(n6592), .S(n5850), .Z(n4372) );
  MUX2_X1 U4969 ( .A(n5362), .B(n6593), .S(n5850), .Z(n4371) );
  MUX2_X1 U4970 ( .A(n5363), .B(n6594), .S(n5850), .Z(n4370) );
  MUX2_X1 U4971 ( .A(n5364), .B(n6595), .S(n5850), .Z(n4369) );
  OAI211_X1 U4972 ( .C1(n6472), .C2(n6621), .A(n6625), .B(n6455), .ZN(n6624)
         );
  NAND3_X1 U4973 ( .A1(n6609), .A2(n6623), .A3(n6610), .ZN(n6625) );
  MUX2_X1 U4974 ( .A(n6531), .B(n5623), .S(n6626), .Z(n4368) );
  MUX2_X1 U4975 ( .A(n6533), .B(n5624), .S(n6626), .Z(n4367) );
  MUX2_X1 U4976 ( .A(n6534), .B(n5625), .S(n6626), .Z(n4366) );
  MUX2_X1 U4977 ( .A(n6535), .B(n5626), .S(n6626), .Z(n4365) );
  MUX2_X1 U4978 ( .A(n6536), .B(n5627), .S(n6626), .Z(n4364) );
  MUX2_X1 U4979 ( .A(n6537), .B(n5628), .S(n6626), .Z(n4363) );
  MUX2_X1 U4980 ( .A(n6538), .B(n5629), .S(n6626), .Z(n4362) );
  MUX2_X1 U4981 ( .A(n6539), .B(n5630), .S(n6626), .Z(n4361) );
  MUX2_X1 U4982 ( .A(n6540), .B(n5631), .S(n6626), .Z(n4360) );
  MUX2_X1 U4983 ( .A(n6541), .B(n5632), .S(n6626), .Z(n4359) );
  MUX2_X1 U4984 ( .A(n6542), .B(n5633), .S(n6626), .Z(n4358) );
  MUX2_X1 U4985 ( .A(n6543), .B(n5634), .S(n6626), .Z(n4357) );
  MUX2_X1 U4986 ( .A(n6544), .B(n5635), .S(n6626), .Z(n4356) );
  MUX2_X1 U4987 ( .A(n6545), .B(n5636), .S(n6626), .Z(n4355) );
  MUX2_X1 U4988 ( .A(n6546), .B(n5637), .S(n6626), .Z(n4354) );
  MUX2_X1 U4989 ( .A(n6547), .B(n5638), .S(n6626), .Z(n4353) );
  MUX2_X1 U4990 ( .A(n6548), .B(n5639), .S(n6626), .Z(n4352) );
  MUX2_X1 U4991 ( .A(n6549), .B(n5640), .S(n6626), .Z(n4351) );
  MUX2_X1 U4992 ( .A(n6550), .B(n5641), .S(n6626), .Z(n4350) );
  MUX2_X1 U4993 ( .A(n6551), .B(n5642), .S(n6626), .Z(n4349) );
  MUX2_X1 U4994 ( .A(n6552), .B(n5643), .S(n6626), .Z(n4348) );
  MUX2_X1 U4995 ( .A(n6553), .B(n5644), .S(n6626), .Z(n4347) );
  MUX2_X1 U4996 ( .A(n6554), .B(n5645), .S(n6626), .Z(n4346) );
  MUX2_X1 U4997 ( .A(n6555), .B(n5646), .S(n6626), .Z(n4345) );
  MUX2_X1 U4998 ( .A(n6556), .B(n5647), .S(n6626), .Z(n4344) );
  MUX2_X1 U4999 ( .A(n6557), .B(n5648), .S(n6626), .Z(n4343) );
  MUX2_X1 U5000 ( .A(n6558), .B(n5649), .S(n6626), .Z(n4342) );
  MUX2_X1 U5001 ( .A(n6559), .B(n5650), .S(n6626), .Z(n4341) );
  MUX2_X1 U5002 ( .A(n6560), .B(n5651), .S(n6626), .Z(n4340) );
  MUX2_X1 U5003 ( .A(n6561), .B(n5652), .S(n6626), .Z(n4339) );
  MUX2_X1 U5004 ( .A(n6562), .B(n5653), .S(n6626), .Z(n4338) );
  MUX2_X1 U5005 ( .A(n6563), .B(n5654), .S(n6626), .Z(n4337) );
  MUX2_X1 U5006 ( .A(n6564), .B(n5655), .S(n6626), .Z(n4336) );
  MUX2_X1 U5007 ( .A(n6565), .B(n5656), .S(n6626), .Z(n4335) );
  MUX2_X1 U5008 ( .A(n6566), .B(n5657), .S(n6626), .Z(n4334) );
  MUX2_X1 U5009 ( .A(n6567), .B(n5658), .S(n6626), .Z(n4333) );
  MUX2_X1 U5010 ( .A(n6568), .B(n5659), .S(n6626), .Z(n4332) );
  MUX2_X1 U5011 ( .A(n6569), .B(n5660), .S(n6626), .Z(n4331) );
  MUX2_X1 U5012 ( .A(n6570), .B(n5661), .S(n6626), .Z(n4330) );
  MUX2_X1 U5013 ( .A(n6571), .B(n5662), .S(n6626), .Z(n4329) );
  MUX2_X1 U5014 ( .A(n6572), .B(n5663), .S(n6626), .Z(n4328) );
  MUX2_X1 U5015 ( .A(n6573), .B(n5664), .S(n6626), .Z(n4327) );
  MUX2_X1 U5016 ( .A(n6574), .B(n5665), .S(n6626), .Z(n4326) );
  MUX2_X1 U5017 ( .A(n6575), .B(n5666), .S(n6626), .Z(n4325) );
  MUX2_X1 U5018 ( .A(n6576), .B(n5667), .S(n6626), .Z(n4324) );
  MUX2_X1 U5019 ( .A(n6577), .B(n5668), .S(n6626), .Z(n4323) );
  MUX2_X1 U5020 ( .A(n6578), .B(n5669), .S(n6626), .Z(n4322) );
  MUX2_X1 U5021 ( .A(n6579), .B(n5670), .S(n6626), .Z(n4321) );
  MUX2_X1 U5022 ( .A(n6580), .B(n5671), .S(n6626), .Z(n4320) );
  MUX2_X1 U5023 ( .A(n6581), .B(n5672), .S(n6626), .Z(n4319) );
  MUX2_X1 U5024 ( .A(n6582), .B(n5673), .S(n6626), .Z(n4318) );
  MUX2_X1 U5025 ( .A(n6583), .B(n5674), .S(n6626), .Z(n4317) );
  MUX2_X1 U5026 ( .A(n6584), .B(n5675), .S(n6626), .Z(n4316) );
  MUX2_X1 U5027 ( .A(n6585), .B(n5676), .S(n6626), .Z(n4315) );
  MUX2_X1 U5028 ( .A(n6586), .B(n5677), .S(n6626), .Z(n4314) );
  MUX2_X1 U5029 ( .A(n6587), .B(n5678), .S(n6626), .Z(n4313) );
  MUX2_X1 U5030 ( .A(n6588), .B(n5679), .S(n6626), .Z(n4312) );
  MUX2_X1 U5031 ( .A(n6589), .B(n5680), .S(n6626), .Z(n4311) );
  MUX2_X1 U5032 ( .A(n6590), .B(n5681), .S(n6626), .Z(n4310) );
  MUX2_X1 U5033 ( .A(n6591), .B(n5682), .S(n6626), .Z(n4309) );
  MUX2_X1 U5034 ( .A(n6592), .B(n5683), .S(n6626), .Z(n4308) );
  MUX2_X1 U5035 ( .A(n6593), .B(n5684), .S(n6626), .Z(n4307) );
  MUX2_X1 U5036 ( .A(n6594), .B(n5685), .S(n6626), .Z(n4306) );
  MUX2_X1 U5037 ( .A(n6595), .B(n5686), .S(n6626), .Z(n4305) );
  AND2_X1 U5038 ( .A1(n6609), .A2(n6629), .ZN(n6605) );
  MUX2_X1 U5039 ( .A(n6531), .B(n8244), .S(n6630), .Z(n4304) );
  MUX2_X1 U5040 ( .A(n6533), .B(n8243), .S(n6630), .Z(n4303) );
  MUX2_X1 U5041 ( .A(n6534), .B(n8242), .S(n6630), .Z(n4302) );
  MUX2_X1 U5042 ( .A(n6535), .B(n8241), .S(n6630), .Z(n4301) );
  MUX2_X1 U5043 ( .A(n6536), .B(n8240), .S(n6630), .Z(n4300) );
  MUX2_X1 U5044 ( .A(n6537), .B(n8239), .S(n6630), .Z(n4299) );
  MUX2_X1 U5045 ( .A(n6538), .B(n8238), .S(n6630), .Z(n4298) );
  MUX2_X1 U5046 ( .A(n6539), .B(n8237), .S(n6630), .Z(n4297) );
  MUX2_X1 U5047 ( .A(n6540), .B(n8236), .S(n6630), .Z(n4296) );
  MUX2_X1 U5048 ( .A(n6541), .B(n8235), .S(n6630), .Z(n4295) );
  MUX2_X1 U5049 ( .A(n6542), .B(n8234), .S(n6630), .Z(n4294) );
  MUX2_X1 U5050 ( .A(n6543), .B(n8233), .S(n6630), .Z(n4293) );
  MUX2_X1 U5051 ( .A(n6544), .B(n8232), .S(n6630), .Z(n4292) );
  MUX2_X1 U5052 ( .A(n6545), .B(n8231), .S(n6630), .Z(n4291) );
  MUX2_X1 U5053 ( .A(n6546), .B(n8230), .S(n6630), .Z(n4290) );
  MUX2_X1 U5054 ( .A(n6547), .B(n8229), .S(n6630), .Z(n4289) );
  MUX2_X1 U5055 ( .A(n6548), .B(n8228), .S(n6630), .Z(n4288) );
  MUX2_X1 U5056 ( .A(n6549), .B(n8227), .S(n6630), .Z(n4287) );
  MUX2_X1 U5057 ( .A(n6550), .B(n8226), .S(n6630), .Z(n4286) );
  MUX2_X1 U5058 ( .A(n6551), .B(n8225), .S(n6630), .Z(n4285) );
  MUX2_X1 U5059 ( .A(n6552), .B(n8224), .S(n6630), .Z(n4284) );
  MUX2_X1 U5060 ( .A(n6553), .B(n8223), .S(n6630), .Z(n4283) );
  MUX2_X1 U5061 ( .A(n6554), .B(n8222), .S(n6630), .Z(n4282) );
  MUX2_X1 U5062 ( .A(n6555), .B(n8221), .S(n6630), .Z(n4281) );
  MUX2_X1 U5063 ( .A(n6556), .B(n8220), .S(n6630), .Z(n4280) );
  MUX2_X1 U5064 ( .A(n6557), .B(n8219), .S(n6630), .Z(n4279) );
  MUX2_X1 U5065 ( .A(n6558), .B(n8218), .S(n6630), .Z(n4278) );
  MUX2_X1 U5066 ( .A(n6559), .B(n8217), .S(n6630), .Z(n4277) );
  MUX2_X1 U5067 ( .A(n6560), .B(n8216), .S(n6630), .Z(n4276) );
  MUX2_X1 U5068 ( .A(n6561), .B(n8215), .S(n6630), .Z(n4275) );
  MUX2_X1 U5069 ( .A(n6562), .B(n8214), .S(n6630), .Z(n4274) );
  MUX2_X1 U5070 ( .A(n6563), .B(n8213), .S(n6630), .Z(n4273) );
  MUX2_X1 U5071 ( .A(n6564), .B(n8212), .S(n6630), .Z(n4272) );
  MUX2_X1 U5072 ( .A(n6565), .B(n8211), .S(n6630), .Z(n4271) );
  MUX2_X1 U5073 ( .A(n6566), .B(n8210), .S(n6630), .Z(n4270) );
  MUX2_X1 U5074 ( .A(n6567), .B(n8209), .S(n6630), .Z(n4269) );
  MUX2_X1 U5075 ( .A(n6568), .B(n8208), .S(n6630), .Z(n4268) );
  MUX2_X1 U5076 ( .A(n6569), .B(n8207), .S(n6630), .Z(n4267) );
  MUX2_X1 U5077 ( .A(n6570), .B(n8206), .S(n6630), .Z(n4266) );
  MUX2_X1 U5078 ( .A(n6571), .B(n8205), .S(n6630), .Z(n4265) );
  MUX2_X1 U5079 ( .A(n6572), .B(n8204), .S(n6630), .Z(n4264) );
  MUX2_X1 U5080 ( .A(n6573), .B(n8203), .S(n6630), .Z(n4263) );
  MUX2_X1 U5081 ( .A(n6574), .B(n8202), .S(n6630), .Z(n4262) );
  MUX2_X1 U5082 ( .A(n6575), .B(n8201), .S(n6630), .Z(n4261) );
  MUX2_X1 U5083 ( .A(n6576), .B(n8200), .S(n6630), .Z(n4260) );
  MUX2_X1 U5084 ( .A(n6577), .B(n8199), .S(n6630), .Z(n4259) );
  MUX2_X1 U5085 ( .A(n6578), .B(n8198), .S(n6630), .Z(n4258) );
  MUX2_X1 U5086 ( .A(n6579), .B(n8197), .S(n6630), .Z(n4257) );
  MUX2_X1 U5087 ( .A(n6580), .B(n8196), .S(n6630), .Z(n4256) );
  MUX2_X1 U5088 ( .A(n6581), .B(n8195), .S(n6630), .Z(n4255) );
  MUX2_X1 U5089 ( .A(n6582), .B(n8194), .S(n6630), .Z(n4254) );
  MUX2_X1 U5090 ( .A(n6583), .B(n8193), .S(n6630), .Z(n4253) );
  MUX2_X1 U5091 ( .A(n6584), .B(n8192), .S(n6630), .Z(n4252) );
  MUX2_X1 U5092 ( .A(n6585), .B(n8191), .S(n6630), .Z(n4251) );
  MUX2_X1 U5093 ( .A(n6586), .B(n8190), .S(n6630), .Z(n4250) );
  MUX2_X1 U5094 ( .A(n6587), .B(n8189), .S(n6630), .Z(n4249) );
  MUX2_X1 U5095 ( .A(n6588), .B(n8188), .S(n6630), .Z(n4248) );
  MUX2_X1 U5096 ( .A(n6589), .B(n8187), .S(n6630), .Z(n4247) );
  MUX2_X1 U5097 ( .A(n6590), .B(n8186), .S(n6630), .Z(n4246) );
  MUX2_X1 U5098 ( .A(n6591), .B(n8185), .S(n6630), .Z(n4245) );
  MUX2_X1 U5099 ( .A(n6592), .B(n8184), .S(n6630), .Z(n4244) );
  MUX2_X1 U5100 ( .A(n6593), .B(n8183), .S(n6630), .Z(n4243) );
  MUX2_X1 U5101 ( .A(n6594), .B(n8182), .S(n6630), .Z(n4242) );
  MUX2_X1 U5102 ( .A(n6595), .B(n8181), .S(n6630), .Z(n4241) );
  INV_X1 U5103 ( .A(n6621), .ZN(n6628) );
  NAND2_X1 U5104 ( .A1(n6617), .A2(n6469), .ZN(n6621) );
  NOR2_X1 U5105 ( .A1(n6618), .A2(N209), .ZN(n6469) );
  INV_X1 U5106 ( .A(N210), .ZN(n6618) );
  NOR2_X1 U5107 ( .A1(n6599), .A2(n6598), .ZN(n6609) );
  INV_X1 U5108 ( .A(n6631), .ZN(n6599) );
  MUX2_X1 U5109 ( .A(n8180), .B(n6531), .S(n5836), .Z(n4240) );
  MUX2_X1 U5110 ( .A(n8179), .B(n6533), .S(n5836), .Z(n4239) );
  MUX2_X1 U5111 ( .A(n8178), .B(n6534), .S(n5836), .Z(n4238) );
  MUX2_X1 U5112 ( .A(n8177), .B(n6535), .S(n5836), .Z(n4237) );
  MUX2_X1 U5113 ( .A(n8176), .B(n6536), .S(n5836), .Z(n4236) );
  MUX2_X1 U5114 ( .A(n8175), .B(n6537), .S(n5836), .Z(n4235) );
  MUX2_X1 U5115 ( .A(n8174), .B(n6538), .S(n5836), .Z(n4234) );
  MUX2_X1 U5116 ( .A(n8173), .B(n6539), .S(n5836), .Z(n4233) );
  MUX2_X1 U5117 ( .A(n8172), .B(n6540), .S(n5836), .Z(n4232) );
  MUX2_X1 U5118 ( .A(n8171), .B(n6541), .S(n5836), .Z(n4231) );
  MUX2_X1 U5119 ( .A(n8170), .B(n6542), .S(n5836), .Z(n4230) );
  MUX2_X1 U5120 ( .A(n8169), .B(n6543), .S(n5836), .Z(n4229) );
  MUX2_X1 U5121 ( .A(n8168), .B(n6544), .S(n5836), .Z(n4228) );
  MUX2_X1 U5122 ( .A(n8167), .B(n6545), .S(n5836), .Z(n4227) );
  MUX2_X1 U5123 ( .A(n8166), .B(n6546), .S(n5836), .Z(n4226) );
  MUX2_X1 U5124 ( .A(n8165), .B(n6547), .S(n5836), .Z(n4225) );
  MUX2_X1 U5125 ( .A(n8164), .B(n6548), .S(n5836), .Z(n4224) );
  MUX2_X1 U5126 ( .A(n8163), .B(n6549), .S(n5836), .Z(n4223) );
  MUX2_X1 U5127 ( .A(n8162), .B(n6550), .S(n5836), .Z(n4222) );
  MUX2_X1 U5128 ( .A(n8161), .B(n6551), .S(n5836), .Z(n4221) );
  MUX2_X1 U5129 ( .A(n8160), .B(n6552), .S(n5836), .Z(n4220) );
  MUX2_X1 U5130 ( .A(n8159), .B(n6553), .S(n5836), .Z(n4219) );
  MUX2_X1 U5131 ( .A(n8158), .B(n6554), .S(n5836), .Z(n4218) );
  MUX2_X1 U5132 ( .A(n8157), .B(n6555), .S(n5836), .Z(n4217) );
  MUX2_X1 U5133 ( .A(n8156), .B(n6556), .S(n5836), .Z(n4216) );
  MUX2_X1 U5134 ( .A(n8155), .B(n6557), .S(n5836), .Z(n4215) );
  MUX2_X1 U5135 ( .A(n8154), .B(n6558), .S(n5836), .Z(n4214) );
  MUX2_X1 U5136 ( .A(n8153), .B(n6559), .S(n5836), .Z(n4213) );
  MUX2_X1 U5137 ( .A(n8152), .B(n6560), .S(n5836), .Z(n4212) );
  MUX2_X1 U5138 ( .A(n8151), .B(n6561), .S(n5836), .Z(n4211) );
  MUX2_X1 U5139 ( .A(n8150), .B(n6562), .S(n5836), .Z(n4210) );
  MUX2_X1 U5140 ( .A(n8149), .B(n6563), .S(n5836), .Z(n4209) );
  MUX2_X1 U5141 ( .A(n8148), .B(n6564), .S(n5836), .Z(n4208) );
  MUX2_X1 U5142 ( .A(n8147), .B(n6565), .S(n5836), .Z(n4207) );
  MUX2_X1 U5143 ( .A(n8146), .B(n6566), .S(n5836), .Z(n4206) );
  MUX2_X1 U5144 ( .A(n8145), .B(n6567), .S(n5836), .Z(n4205) );
  MUX2_X1 U5145 ( .A(n8144), .B(n6568), .S(n5836), .Z(n4204) );
  MUX2_X1 U5146 ( .A(n8143), .B(n6569), .S(n5836), .Z(n4203) );
  MUX2_X1 U5147 ( .A(n8142), .B(n6570), .S(n5836), .Z(n4202) );
  MUX2_X1 U5148 ( .A(n8141), .B(n6571), .S(n5836), .Z(n4201) );
  MUX2_X1 U5149 ( .A(n8140), .B(n6572), .S(n5836), .Z(n4200) );
  MUX2_X1 U5150 ( .A(n8139), .B(n6573), .S(n5836), .Z(n4199) );
  MUX2_X1 U5151 ( .A(n8138), .B(n6574), .S(n5836), .Z(n4198) );
  MUX2_X1 U5152 ( .A(n8137), .B(n6575), .S(n5836), .Z(n4197) );
  MUX2_X1 U5153 ( .A(n8136), .B(n6576), .S(n5836), .Z(n4196) );
  MUX2_X1 U5154 ( .A(n8135), .B(n6577), .S(n5836), .Z(n4195) );
  MUX2_X1 U5155 ( .A(n8134), .B(n6578), .S(n5836), .Z(n4194) );
  MUX2_X1 U5156 ( .A(n8133), .B(n6579), .S(n5836), .Z(n4193) );
  MUX2_X1 U5157 ( .A(n8132), .B(n6580), .S(n5836), .Z(n4192) );
  MUX2_X1 U5158 ( .A(n8131), .B(n6581), .S(n5836), .Z(n4191) );
  MUX2_X1 U5159 ( .A(n8130), .B(n6582), .S(n5836), .Z(n4190) );
  MUX2_X1 U5160 ( .A(n8129), .B(n6583), .S(n5836), .Z(n4189) );
  MUX2_X1 U5161 ( .A(n8128), .B(n6584), .S(n5836), .Z(n4188) );
  MUX2_X1 U5162 ( .A(n8127), .B(n6585), .S(n5836), .Z(n4187) );
  MUX2_X1 U5163 ( .A(n8126), .B(n6586), .S(n5836), .Z(n4186) );
  MUX2_X1 U5164 ( .A(n8125), .B(n6587), .S(n5836), .Z(n4185) );
  MUX2_X1 U5165 ( .A(n8124), .B(n6588), .S(n5836), .Z(n4184) );
  MUX2_X1 U5166 ( .A(n8123), .B(n6589), .S(n5836), .Z(n4183) );
  MUX2_X1 U5167 ( .A(n8122), .B(n6590), .S(n5836), .Z(n4182) );
  MUX2_X1 U5168 ( .A(n8121), .B(n6591), .S(n5836), .Z(n4181) );
  MUX2_X1 U5169 ( .A(n8120), .B(n6592), .S(n5836), .Z(n4180) );
  MUX2_X1 U5170 ( .A(n8119), .B(n6593), .S(n5836), .Z(n4179) );
  MUX2_X1 U5171 ( .A(n8118), .B(n6594), .S(n5836), .Z(n4178) );
  MUX2_X1 U5172 ( .A(n8117), .B(n6595), .S(n5836), .Z(n4177) );
  OAI211_X1 U5173 ( .C1(n6473), .C2(n6633), .A(n6634), .B(n6455), .ZN(n6632)
         );
  NAND3_X1 U5174 ( .A1(n6604), .A2(n6606), .A3(n6635), .ZN(n6634) );
  MUX2_X1 U5175 ( .A(n5751), .B(n6531), .S(n5838), .Z(n4176) );
  MUX2_X1 U5176 ( .A(n5752), .B(n6533), .S(n5838), .Z(n4175) );
  MUX2_X1 U5177 ( .A(n5753), .B(n6534), .S(n5838), .Z(n4174) );
  MUX2_X1 U5178 ( .A(n5754), .B(n6535), .S(n5838), .Z(n4173) );
  MUX2_X1 U5179 ( .A(n5755), .B(n6536), .S(n5838), .Z(n4172) );
  MUX2_X1 U5180 ( .A(n5756), .B(n6537), .S(n5838), .Z(n4171) );
  MUX2_X1 U5181 ( .A(n5757), .B(n6538), .S(n5838), .Z(n4170) );
  MUX2_X1 U5182 ( .A(n5758), .B(n6539), .S(n5838), .Z(n4169) );
  MUX2_X1 U5183 ( .A(n5759), .B(n6540), .S(n5838), .Z(n4168) );
  MUX2_X1 U5184 ( .A(n5760), .B(n6541), .S(n5838), .Z(n4167) );
  MUX2_X1 U5185 ( .A(n5761), .B(n6542), .S(n5838), .Z(n4166) );
  MUX2_X1 U5186 ( .A(n5762), .B(n6543), .S(n5838), .Z(n4165) );
  MUX2_X1 U5187 ( .A(n5763), .B(n6544), .S(n5838), .Z(n4164) );
  MUX2_X1 U5188 ( .A(n5764), .B(n6545), .S(n5838), .Z(n4163) );
  MUX2_X1 U5189 ( .A(n5765), .B(n6546), .S(n5838), .Z(n4162) );
  MUX2_X1 U5190 ( .A(n5766), .B(n6547), .S(n5838), .Z(n4161) );
  MUX2_X1 U5191 ( .A(n5767), .B(n6548), .S(n5838), .Z(n4160) );
  MUX2_X1 U5192 ( .A(n5768), .B(n6549), .S(n5838), .Z(n4159) );
  MUX2_X1 U5193 ( .A(n5769), .B(n6550), .S(n5838), .Z(n4158) );
  MUX2_X1 U5194 ( .A(n5770), .B(n6551), .S(n5838), .Z(n4157) );
  MUX2_X1 U5195 ( .A(n5771), .B(n6552), .S(n5838), .Z(n4156) );
  MUX2_X1 U5196 ( .A(n5772), .B(n6553), .S(n5838), .Z(n4155) );
  MUX2_X1 U5197 ( .A(n5773), .B(n6554), .S(n5838), .Z(n4154) );
  MUX2_X1 U5198 ( .A(n5774), .B(n6555), .S(n5838), .Z(n4153) );
  MUX2_X1 U5199 ( .A(n5775), .B(n6556), .S(n5838), .Z(n4152) );
  MUX2_X1 U5200 ( .A(n5776), .B(n6557), .S(n5838), .Z(n4151) );
  MUX2_X1 U5201 ( .A(n5777), .B(n6558), .S(n5838), .Z(n4150) );
  MUX2_X1 U5202 ( .A(n5778), .B(n6559), .S(n5838), .Z(n4149) );
  MUX2_X1 U5203 ( .A(n5779), .B(n6560), .S(n5838), .Z(n4148) );
  MUX2_X1 U5204 ( .A(n5780), .B(n6561), .S(n5838), .Z(n4147) );
  MUX2_X1 U5205 ( .A(n5781), .B(n6562), .S(n5838), .Z(n4146) );
  MUX2_X1 U5206 ( .A(n5782), .B(n6563), .S(n5838), .Z(n4145) );
  MUX2_X1 U5207 ( .A(n5783), .B(n6564), .S(n5838), .Z(n4144) );
  MUX2_X1 U5208 ( .A(n5784), .B(n6565), .S(n5838), .Z(n4143) );
  MUX2_X1 U5209 ( .A(n5785), .B(n6566), .S(n5838), .Z(n4142) );
  MUX2_X1 U5210 ( .A(n5786), .B(n6567), .S(n5838), .Z(n4141) );
  MUX2_X1 U5211 ( .A(n5787), .B(n6568), .S(n5838), .Z(n4140) );
  MUX2_X1 U5212 ( .A(n5788), .B(n6569), .S(n5838), .Z(n4139) );
  MUX2_X1 U5213 ( .A(n5789), .B(n6570), .S(n5838), .Z(n4138) );
  MUX2_X1 U5214 ( .A(n5790), .B(n6571), .S(n5838), .Z(n4137) );
  MUX2_X1 U5215 ( .A(n5791), .B(n6572), .S(n5838), .Z(n4136) );
  MUX2_X1 U5216 ( .A(n5792), .B(n6573), .S(n5838), .Z(n4135) );
  MUX2_X1 U5217 ( .A(n5793), .B(n6574), .S(n5838), .Z(n4134) );
  MUX2_X1 U5218 ( .A(n5794), .B(n6575), .S(n5838), .Z(n4133) );
  MUX2_X1 U5219 ( .A(n5795), .B(n6576), .S(n5838), .Z(n4132) );
  MUX2_X1 U5220 ( .A(n5796), .B(n6577), .S(n5838), .Z(n4131) );
  MUX2_X1 U5221 ( .A(n5797), .B(n6578), .S(n5838), .Z(n4130) );
  MUX2_X1 U5222 ( .A(n5798), .B(n6579), .S(n5838), .Z(n4129) );
  MUX2_X1 U5223 ( .A(n5799), .B(n6580), .S(n5838), .Z(n4128) );
  MUX2_X1 U5224 ( .A(n5800), .B(n6581), .S(n5838), .Z(n4127) );
  MUX2_X1 U5225 ( .A(n5801), .B(n6582), .S(n5838), .Z(n4126) );
  MUX2_X1 U5226 ( .A(n5802), .B(n6583), .S(n5838), .Z(n4125) );
  MUX2_X1 U5227 ( .A(n5803), .B(n6584), .S(n5838), .Z(n4124) );
  MUX2_X1 U5228 ( .A(n5804), .B(n6585), .S(n5838), .Z(n4123) );
  MUX2_X1 U5229 ( .A(n5805), .B(n6586), .S(n5838), .Z(n4122) );
  MUX2_X1 U5230 ( .A(n5806), .B(n6587), .S(n5838), .Z(n4121) );
  MUX2_X1 U5231 ( .A(n5807), .B(n6588), .S(n5838), .Z(n4120) );
  MUX2_X1 U5232 ( .A(n5808), .B(n6589), .S(n5838), .Z(n4119) );
  MUX2_X1 U5233 ( .A(n5809), .B(n6590), .S(n5838), .Z(n4118) );
  MUX2_X1 U5234 ( .A(n5810), .B(n6591), .S(n5838), .Z(n4117) );
  MUX2_X1 U5235 ( .A(n5811), .B(n6592), .S(n5838), .Z(n4116) );
  MUX2_X1 U5236 ( .A(n5812), .B(n6593), .S(n5838), .Z(n4115) );
  MUX2_X1 U5237 ( .A(n5813), .B(n6594), .S(n5838), .Z(n4114) );
  MUX2_X1 U5238 ( .A(n5814), .B(n6595), .S(n5838), .Z(n4113) );
  OAI211_X1 U5239 ( .C1(n6472), .C2(n6633), .A(n6637), .B(n6455), .ZN(n6636)
         );
  NAND3_X1 U5240 ( .A1(n6610), .A2(n6606), .A3(n6638), .ZN(n6637) );
  MUX2_X1 U5241 ( .A(n6531), .B(n5559), .S(n6639), .Z(n4112) );
  MUX2_X1 U5242 ( .A(n6533), .B(n5560), .S(n6639), .Z(n4111) );
  MUX2_X1 U5243 ( .A(n6534), .B(n5561), .S(n6639), .Z(n4110) );
  MUX2_X1 U5244 ( .A(n6535), .B(n5562), .S(n6639), .Z(n4109) );
  MUX2_X1 U5245 ( .A(n6536), .B(n5563), .S(n6639), .Z(n4108) );
  MUX2_X1 U5246 ( .A(n6537), .B(n5564), .S(n6639), .Z(n4107) );
  MUX2_X1 U5247 ( .A(n6538), .B(n5565), .S(n6639), .Z(n4106) );
  MUX2_X1 U5248 ( .A(n6539), .B(n5566), .S(n6639), .Z(n4105) );
  MUX2_X1 U5249 ( .A(n6540), .B(n5567), .S(n6639), .Z(n4104) );
  MUX2_X1 U5250 ( .A(n6541), .B(n5568), .S(n6639), .Z(n4103) );
  MUX2_X1 U5251 ( .A(n6542), .B(n5569), .S(n6639), .Z(n4102) );
  MUX2_X1 U5252 ( .A(n6543), .B(n5570), .S(n6639), .Z(n4101) );
  MUX2_X1 U5253 ( .A(n6544), .B(n5571), .S(n6639), .Z(n4100) );
  MUX2_X1 U5254 ( .A(n6545), .B(n5572), .S(n6639), .Z(n4099) );
  MUX2_X1 U5255 ( .A(n6546), .B(n5573), .S(n6639), .Z(n4098) );
  MUX2_X1 U5256 ( .A(n6547), .B(n5574), .S(n6639), .Z(n4097) );
  MUX2_X1 U5257 ( .A(n6548), .B(n5575), .S(n6639), .Z(n4096) );
  MUX2_X1 U5258 ( .A(n6549), .B(n5576), .S(n6639), .Z(n4095) );
  MUX2_X1 U5259 ( .A(n6550), .B(n5577), .S(n6639), .Z(n4094) );
  MUX2_X1 U5260 ( .A(n6551), .B(n5578), .S(n6639), .Z(n4093) );
  MUX2_X1 U5261 ( .A(n6552), .B(n5579), .S(n6639), .Z(n4092) );
  MUX2_X1 U5262 ( .A(n6553), .B(n5580), .S(n6639), .Z(n4091) );
  MUX2_X1 U5263 ( .A(n6554), .B(n5581), .S(n6639), .Z(n4090) );
  MUX2_X1 U5264 ( .A(n6555), .B(n5582), .S(n6639), .Z(n4089) );
  MUX2_X1 U5265 ( .A(n6556), .B(n5583), .S(n6639), .Z(n4088) );
  MUX2_X1 U5266 ( .A(n6557), .B(n5584), .S(n6639), .Z(n4087) );
  MUX2_X1 U5267 ( .A(n6558), .B(n5585), .S(n6639), .Z(n4086) );
  MUX2_X1 U5268 ( .A(n6559), .B(n5586), .S(n6639), .Z(n4085) );
  MUX2_X1 U5269 ( .A(n6560), .B(n5587), .S(n6639), .Z(n4084) );
  MUX2_X1 U5270 ( .A(n6561), .B(n5588), .S(n6639), .Z(n4083) );
  MUX2_X1 U5271 ( .A(n6562), .B(n5589), .S(n6639), .Z(n4082) );
  MUX2_X1 U5272 ( .A(n6563), .B(n5590), .S(n6639), .Z(n4081) );
  MUX2_X1 U5273 ( .A(n6564), .B(n5591), .S(n6639), .Z(n4080) );
  MUX2_X1 U5274 ( .A(n6565), .B(n5592), .S(n6639), .Z(n4079) );
  MUX2_X1 U5275 ( .A(n6566), .B(n5593), .S(n6639), .Z(n4078) );
  MUX2_X1 U5276 ( .A(n6567), .B(n5594), .S(n6639), .Z(n4077) );
  MUX2_X1 U5277 ( .A(n6568), .B(n5595), .S(n6639), .Z(n4076) );
  MUX2_X1 U5278 ( .A(n6569), .B(n5596), .S(n6639), .Z(n4075) );
  MUX2_X1 U5279 ( .A(n6570), .B(n5597), .S(n6639), .Z(n4074) );
  MUX2_X1 U5280 ( .A(n6571), .B(n5598), .S(n6639), .Z(n4073) );
  MUX2_X1 U5281 ( .A(n6572), .B(n5599), .S(n6639), .Z(n4072) );
  MUX2_X1 U5282 ( .A(n6573), .B(n5600), .S(n6639), .Z(n4071) );
  MUX2_X1 U5283 ( .A(n6574), .B(n5601), .S(n6639), .Z(n4070) );
  MUX2_X1 U5284 ( .A(n6575), .B(n5602), .S(n6639), .Z(n4069) );
  MUX2_X1 U5285 ( .A(n6576), .B(n5603), .S(n6639), .Z(n4068) );
  MUX2_X1 U5286 ( .A(n6577), .B(n5604), .S(n6639), .Z(n4067) );
  MUX2_X1 U5287 ( .A(n6578), .B(n5605), .S(n6639), .Z(n4066) );
  MUX2_X1 U5288 ( .A(n6579), .B(n5606), .S(n6639), .Z(n4065) );
  MUX2_X1 U5289 ( .A(n6580), .B(n5607), .S(n6639), .Z(n4064) );
  MUX2_X1 U5290 ( .A(n6581), .B(n5608), .S(n6639), .Z(n4063) );
  MUX2_X1 U5291 ( .A(n6582), .B(n5609), .S(n6639), .Z(n4062) );
  MUX2_X1 U5292 ( .A(n6583), .B(n5610), .S(n6639), .Z(n4061) );
  MUX2_X1 U5293 ( .A(n6584), .B(n5611), .S(n6639), .Z(n4060) );
  MUX2_X1 U5294 ( .A(n6585), .B(n5612), .S(n6639), .Z(n4059) );
  MUX2_X1 U5295 ( .A(n6586), .B(n5613), .S(n6639), .Z(n4058) );
  MUX2_X1 U5296 ( .A(n6587), .B(n5614), .S(n6639), .Z(n4057) );
  MUX2_X1 U5297 ( .A(n6588), .B(n5615), .S(n6639), .Z(n4056) );
  MUX2_X1 U5298 ( .A(n6589), .B(n5616), .S(n6639), .Z(n4055) );
  MUX2_X1 U5299 ( .A(n6590), .B(n5617), .S(n6639), .Z(n4054) );
  MUX2_X1 U5300 ( .A(n6591), .B(n5618), .S(n6639), .Z(n4053) );
  MUX2_X1 U5301 ( .A(n6592), .B(n5619), .S(n6639), .Z(n4052) );
  MUX2_X1 U5302 ( .A(n6593), .B(n5620), .S(n6639), .Z(n4051) );
  MUX2_X1 U5303 ( .A(n6594), .B(n5621), .S(n6639), .Z(n4050) );
  MUX2_X1 U5304 ( .A(n6595), .B(n5622), .S(n6639), .Z(n4049) );
  MUX2_X1 U5305 ( .A(n6531), .B(n8116), .S(n6641), .Z(n4048) );
  MUX2_X1 U5306 ( .A(n6533), .B(n8115), .S(n6641), .Z(n4047) );
  MUX2_X1 U5307 ( .A(n6534), .B(n8114), .S(n6641), .Z(n4046) );
  MUX2_X1 U5308 ( .A(n6535), .B(n8113), .S(n6641), .Z(n4045) );
  MUX2_X1 U5309 ( .A(n6536), .B(n8112), .S(n6641), .Z(n4044) );
  MUX2_X1 U5310 ( .A(n6537), .B(n8111), .S(n6641), .Z(n4043) );
  MUX2_X1 U5311 ( .A(n6538), .B(n8110), .S(n6641), .Z(n4042) );
  MUX2_X1 U5312 ( .A(n6539), .B(n8109), .S(n6641), .Z(n4041) );
  MUX2_X1 U5313 ( .A(n6540), .B(n8108), .S(n6641), .Z(n4040) );
  MUX2_X1 U5314 ( .A(n6541), .B(n8107), .S(n6641), .Z(n4039) );
  MUX2_X1 U5315 ( .A(n6542), .B(n8106), .S(n6641), .Z(n4038) );
  MUX2_X1 U5316 ( .A(n6543), .B(n8105), .S(n6641), .Z(n4037) );
  MUX2_X1 U5317 ( .A(n6544), .B(n8104), .S(n6641), .Z(n4036) );
  MUX2_X1 U5318 ( .A(n6545), .B(n8103), .S(n6641), .Z(n4035) );
  MUX2_X1 U5319 ( .A(n6546), .B(n8102), .S(n6641), .Z(n4034) );
  MUX2_X1 U5320 ( .A(n6547), .B(n8101), .S(n6641), .Z(n4033) );
  MUX2_X1 U5321 ( .A(n6548), .B(n8100), .S(n6641), .Z(n4032) );
  MUX2_X1 U5322 ( .A(n6549), .B(n8099), .S(n6641), .Z(n4031) );
  MUX2_X1 U5323 ( .A(n6550), .B(n8098), .S(n6641), .Z(n4030) );
  MUX2_X1 U5324 ( .A(n6551), .B(n8097), .S(n6641), .Z(n4029) );
  MUX2_X1 U5325 ( .A(n6552), .B(n8096), .S(n6641), .Z(n4028) );
  MUX2_X1 U5326 ( .A(n6553), .B(n8095), .S(n6641), .Z(n4027) );
  MUX2_X1 U5327 ( .A(n6554), .B(n8094), .S(n6641), .Z(n4026) );
  MUX2_X1 U5328 ( .A(n6555), .B(n8093), .S(n6641), .Z(n4025) );
  MUX2_X1 U5329 ( .A(n6556), .B(n8092), .S(n6641), .Z(n4024) );
  MUX2_X1 U5330 ( .A(n6557), .B(n8091), .S(n6641), .Z(n4023) );
  MUX2_X1 U5331 ( .A(n6558), .B(n8090), .S(n6641), .Z(n4022) );
  MUX2_X1 U5332 ( .A(n6559), .B(n8089), .S(n6641), .Z(n4021) );
  MUX2_X1 U5333 ( .A(n6560), .B(n8088), .S(n6641), .Z(n4020) );
  MUX2_X1 U5334 ( .A(n6561), .B(n8087), .S(n6641), .Z(n4019) );
  MUX2_X1 U5335 ( .A(n6562), .B(n8086), .S(n6641), .Z(n4018) );
  MUX2_X1 U5336 ( .A(n6563), .B(n8085), .S(n6641), .Z(n4017) );
  MUX2_X1 U5337 ( .A(n6564), .B(n8084), .S(n6641), .Z(n4016) );
  MUX2_X1 U5338 ( .A(n6565), .B(n8083), .S(n6641), .Z(n4015) );
  MUX2_X1 U5339 ( .A(n6566), .B(n8082), .S(n6641), .Z(n4014) );
  MUX2_X1 U5340 ( .A(n6567), .B(n8081), .S(n6641), .Z(n4013) );
  MUX2_X1 U5341 ( .A(n6568), .B(n8080), .S(n6641), .Z(n4012) );
  MUX2_X1 U5342 ( .A(n6569), .B(n8079), .S(n6641), .Z(n4011) );
  MUX2_X1 U5343 ( .A(n6570), .B(n8078), .S(n6641), .Z(n4010) );
  MUX2_X1 U5344 ( .A(n6571), .B(n8077), .S(n6641), .Z(n4009) );
  MUX2_X1 U5345 ( .A(n6572), .B(n8076), .S(n6641), .Z(n4008) );
  MUX2_X1 U5346 ( .A(n6573), .B(n8075), .S(n6641), .Z(n4007) );
  MUX2_X1 U5347 ( .A(n6574), .B(n8074), .S(n6641), .Z(n4006) );
  MUX2_X1 U5348 ( .A(n6575), .B(n8073), .S(n6641), .Z(n4005) );
  MUX2_X1 U5349 ( .A(n6576), .B(n8072), .S(n6641), .Z(n4004) );
  MUX2_X1 U5350 ( .A(n6577), .B(n8071), .S(n6641), .Z(n4003) );
  MUX2_X1 U5351 ( .A(n6578), .B(n8070), .S(n6641), .Z(n4002) );
  MUX2_X1 U5352 ( .A(n6579), .B(n8069), .S(n6641), .Z(n4001) );
  MUX2_X1 U5353 ( .A(n6580), .B(n8068), .S(n6641), .Z(n4000) );
  MUX2_X1 U5354 ( .A(n6581), .B(n8067), .S(n6641), .Z(n3999) );
  MUX2_X1 U5355 ( .A(n6582), .B(n8066), .S(n6641), .Z(n3998) );
  MUX2_X1 U5356 ( .A(n6583), .B(n8065), .S(n6641), .Z(n3997) );
  MUX2_X1 U5357 ( .A(n6584), .B(n8064), .S(n6641), .Z(n3996) );
  MUX2_X1 U5358 ( .A(n6585), .B(n8063), .S(n6641), .Z(n3995) );
  MUX2_X1 U5359 ( .A(n6586), .B(n8062), .S(n6641), .Z(n3994) );
  MUX2_X1 U5360 ( .A(n6587), .B(n8061), .S(n6641), .Z(n3993) );
  MUX2_X1 U5361 ( .A(n6588), .B(n8060), .S(n6641), .Z(n3992) );
  MUX2_X1 U5362 ( .A(n6589), .B(n8059), .S(n6641), .Z(n3991) );
  MUX2_X1 U5363 ( .A(n6590), .B(n8058), .S(n6641), .Z(n3990) );
  MUX2_X1 U5364 ( .A(n6591), .B(n8057), .S(n6641), .Z(n3989) );
  MUX2_X1 U5365 ( .A(n6592), .B(n8056), .S(n6641), .Z(n3988) );
  MUX2_X1 U5366 ( .A(n6593), .B(n8055), .S(n6641), .Z(n3987) );
  MUX2_X1 U5367 ( .A(n6594), .B(n8054), .S(n6641), .Z(n3986) );
  MUX2_X1 U5368 ( .A(n6595), .B(n8053), .S(n6641), .Z(n3985) );
  AND3_X1 U5369 ( .A1(n6612), .A2(n6616), .A3(n6638), .ZN(n6642) );
  AND2_X1 U5370 ( .A1(n6606), .A2(n6643), .ZN(n6612) );
  AND2_X1 U5371 ( .A1(n6644), .A2(n6645), .ZN(n6606) );
  INV_X1 U5372 ( .A(n6633), .ZN(n6640) );
  NAND2_X1 U5373 ( .A1(n6617), .A2(n6466), .ZN(n6633) );
  NOR2_X1 U5374 ( .A1(n6619), .A2(N210), .ZN(n6466) );
  MUX2_X1 U5375 ( .A(n8052), .B(n6531), .S(n5840), .Z(n3984) );
  MUX2_X1 U5376 ( .A(n8051), .B(n6533), .S(n5840), .Z(n3983) );
  MUX2_X1 U5377 ( .A(n8050), .B(n6534), .S(n5840), .Z(n3982) );
  MUX2_X1 U5378 ( .A(n8049), .B(n6535), .S(n5840), .Z(n3981) );
  MUX2_X1 U5379 ( .A(n8048), .B(n6536), .S(n5840), .Z(n3980) );
  MUX2_X1 U5380 ( .A(n8047), .B(n6537), .S(n5840), .Z(n3979) );
  MUX2_X1 U5381 ( .A(n8046), .B(n6538), .S(n5840), .Z(n3978) );
  MUX2_X1 U5382 ( .A(n8045), .B(n6539), .S(n5840), .Z(n3977) );
  MUX2_X1 U5383 ( .A(n8044), .B(n6540), .S(n5840), .Z(n3976) );
  MUX2_X1 U5384 ( .A(n8043), .B(n6541), .S(n5840), .Z(n3975) );
  MUX2_X1 U5385 ( .A(n8042), .B(n6542), .S(n5840), .Z(n3974) );
  MUX2_X1 U5386 ( .A(n8041), .B(n6543), .S(n5840), .Z(n3973) );
  MUX2_X1 U5387 ( .A(n8040), .B(n6544), .S(n5840), .Z(n3972) );
  MUX2_X1 U5388 ( .A(n8039), .B(n6545), .S(n5840), .Z(n3971) );
  MUX2_X1 U5389 ( .A(n8038), .B(n6546), .S(n5840), .Z(n3970) );
  MUX2_X1 U5390 ( .A(n8037), .B(n6547), .S(n5840), .Z(n3969) );
  MUX2_X1 U5391 ( .A(n8036), .B(n6548), .S(n5840), .Z(n3968) );
  MUX2_X1 U5392 ( .A(n8035), .B(n6549), .S(n5840), .Z(n3967) );
  MUX2_X1 U5393 ( .A(n8034), .B(n6550), .S(n5840), .Z(n3966) );
  MUX2_X1 U5394 ( .A(n8033), .B(n6551), .S(n5840), .Z(n3965) );
  MUX2_X1 U5395 ( .A(n8032), .B(n6552), .S(n5840), .Z(n3964) );
  MUX2_X1 U5396 ( .A(n8031), .B(n6553), .S(n5840), .Z(n3963) );
  MUX2_X1 U5397 ( .A(n8030), .B(n6554), .S(n5840), .Z(n3962) );
  MUX2_X1 U5398 ( .A(n8029), .B(n6555), .S(n5840), .Z(n3961) );
  MUX2_X1 U5399 ( .A(n8028), .B(n6556), .S(n5840), .Z(n3960) );
  MUX2_X1 U5400 ( .A(n8027), .B(n6557), .S(n5840), .Z(n3959) );
  MUX2_X1 U5401 ( .A(n8026), .B(n6558), .S(n5840), .Z(n3958) );
  MUX2_X1 U5402 ( .A(n8025), .B(n6559), .S(n5840), .Z(n3957) );
  MUX2_X1 U5403 ( .A(n8024), .B(n6560), .S(n5840), .Z(n3956) );
  MUX2_X1 U5404 ( .A(n8023), .B(n6561), .S(n5840), .Z(n3955) );
  MUX2_X1 U5405 ( .A(n8022), .B(n6562), .S(n5840), .Z(n3954) );
  MUX2_X1 U5406 ( .A(n8021), .B(n6563), .S(n5840), .Z(n3953) );
  MUX2_X1 U5407 ( .A(n8020), .B(n6564), .S(n5840), .Z(n3952) );
  MUX2_X1 U5408 ( .A(n8019), .B(n6565), .S(n5840), .Z(n3951) );
  MUX2_X1 U5409 ( .A(n8018), .B(n6566), .S(n5840), .Z(n3950) );
  MUX2_X1 U5410 ( .A(n8017), .B(n6567), .S(n5840), .Z(n3949) );
  MUX2_X1 U5411 ( .A(n8016), .B(n6568), .S(n5840), .Z(n3948) );
  MUX2_X1 U5412 ( .A(n8015), .B(n6569), .S(n5840), .Z(n3947) );
  MUX2_X1 U5413 ( .A(n8014), .B(n6570), .S(n5840), .Z(n3946) );
  MUX2_X1 U5414 ( .A(n8013), .B(n6571), .S(n5840), .Z(n3945) );
  MUX2_X1 U5415 ( .A(n8012), .B(n6572), .S(n5840), .Z(n3944) );
  MUX2_X1 U5416 ( .A(n8011), .B(n6573), .S(n5840), .Z(n3943) );
  MUX2_X1 U5417 ( .A(n8010), .B(n6574), .S(n5840), .Z(n3942) );
  MUX2_X1 U5418 ( .A(n8009), .B(n6575), .S(n5840), .Z(n3941) );
  MUX2_X1 U5419 ( .A(n8008), .B(n6576), .S(n5840), .Z(n3940) );
  MUX2_X1 U5420 ( .A(n8007), .B(n6577), .S(n5840), .Z(n3939) );
  MUX2_X1 U5421 ( .A(n8006), .B(n6578), .S(n5840), .Z(n3938) );
  MUX2_X1 U5422 ( .A(n8005), .B(n6579), .S(n5840), .Z(n3937) );
  MUX2_X1 U5423 ( .A(n8004), .B(n6580), .S(n5840), .Z(n3936) );
  MUX2_X1 U5424 ( .A(n8003), .B(n6581), .S(n5840), .Z(n3935) );
  MUX2_X1 U5425 ( .A(n8002), .B(n6582), .S(n5840), .Z(n3934) );
  MUX2_X1 U5426 ( .A(n8001), .B(n6583), .S(n5840), .Z(n3933) );
  MUX2_X1 U5427 ( .A(n8000), .B(n6584), .S(n5840), .Z(n3932) );
  MUX2_X1 U5428 ( .A(n7999), .B(n6585), .S(n5840), .Z(n3931) );
  MUX2_X1 U5429 ( .A(n7998), .B(n6586), .S(n5840), .Z(n3930) );
  MUX2_X1 U5430 ( .A(n7997), .B(n6587), .S(n5840), .Z(n3929) );
  MUX2_X1 U5431 ( .A(n7996), .B(n6588), .S(n5840), .Z(n3928) );
  MUX2_X1 U5432 ( .A(n7995), .B(n6589), .S(n5840), .Z(n3927) );
  MUX2_X1 U5433 ( .A(n7994), .B(n6590), .S(n5840), .Z(n3926) );
  MUX2_X1 U5434 ( .A(n7993), .B(n6591), .S(n5840), .Z(n3925) );
  MUX2_X1 U5435 ( .A(n7992), .B(n6592), .S(n5840), .Z(n3924) );
  MUX2_X1 U5436 ( .A(n7991), .B(n6593), .S(n5840), .Z(n3923) );
  MUX2_X1 U5437 ( .A(n7990), .B(n6594), .S(n5840), .Z(n3922) );
  MUX2_X1 U5438 ( .A(n7989), .B(n6595), .S(n5840), .Z(n3921) );
  OAI211_X1 U5439 ( .C1(n6473), .C2(n6647), .A(n6648), .B(n6455), .ZN(n6646)
         );
  NAND3_X1 U5440 ( .A1(n6604), .A2(n6623), .A3(n6635), .ZN(n6648) );
  NAND2_X1 U5441 ( .A1(N208), .A2(n5855), .ZN(n6473) );
  MUX2_X1 U5442 ( .A(n4961), .B(n6531), .S(n5842), .Z(n3920) );
  MUX2_X1 U5443 ( .A(n4962), .B(n6533), .S(n5842), .Z(n3919) );
  MUX2_X1 U5444 ( .A(n4963), .B(n6534), .S(n5842), .Z(n3918) );
  MUX2_X1 U5445 ( .A(n4964), .B(n6535), .S(n5842), .Z(n3917) );
  MUX2_X1 U5446 ( .A(n4965), .B(n6536), .S(n5842), .Z(n3916) );
  MUX2_X1 U5447 ( .A(n4966), .B(n6537), .S(n5842), .Z(n3915) );
  MUX2_X1 U5448 ( .A(n4967), .B(n6538), .S(n5842), .Z(n3914) );
  MUX2_X1 U5449 ( .A(n4968), .B(n6539), .S(n5842), .Z(n3913) );
  MUX2_X1 U5450 ( .A(n4969), .B(n6540), .S(n5842), .Z(n3912) );
  MUX2_X1 U5451 ( .A(n4970), .B(n6541), .S(n5842), .Z(n3911) );
  MUX2_X1 U5452 ( .A(n4971), .B(n6542), .S(n5842), .Z(n3910) );
  MUX2_X1 U5453 ( .A(n4972), .B(n6543), .S(n5842), .Z(n3909) );
  MUX2_X1 U5454 ( .A(n4973), .B(n6544), .S(n5842), .Z(n3908) );
  MUX2_X1 U5455 ( .A(n4974), .B(n6545), .S(n5842), .Z(n3907) );
  MUX2_X1 U5456 ( .A(n4975), .B(n6546), .S(n5842), .Z(n3906) );
  MUX2_X1 U5457 ( .A(n4976), .B(n6547), .S(n5842), .Z(n3905) );
  MUX2_X1 U5458 ( .A(n4977), .B(n6548), .S(n5842), .Z(n3904) );
  MUX2_X1 U5459 ( .A(n4978), .B(n6549), .S(n5842), .Z(n3903) );
  MUX2_X1 U5460 ( .A(n4979), .B(n6550), .S(n5842), .Z(n3902) );
  MUX2_X1 U5461 ( .A(n4980), .B(n6551), .S(n5842), .Z(n3901) );
  MUX2_X1 U5462 ( .A(n4981), .B(n6552), .S(n5842), .Z(n3900) );
  MUX2_X1 U5463 ( .A(n4982), .B(n6553), .S(n5842), .Z(n3899) );
  MUX2_X1 U5464 ( .A(n4983), .B(n6554), .S(n5842), .Z(n3898) );
  MUX2_X1 U5465 ( .A(n4984), .B(n6555), .S(n5842), .Z(n3897) );
  MUX2_X1 U5466 ( .A(n4985), .B(n6556), .S(n5842), .Z(n3896) );
  MUX2_X1 U5467 ( .A(n4986), .B(n6557), .S(n5842), .Z(n3895) );
  MUX2_X1 U5468 ( .A(n4987), .B(n6558), .S(n5842), .Z(n3894) );
  MUX2_X1 U5469 ( .A(n4988), .B(n6559), .S(n5842), .Z(n3893) );
  MUX2_X1 U5470 ( .A(n4989), .B(n6560), .S(n5842), .Z(n3892) );
  MUX2_X1 U5471 ( .A(n4990), .B(n6561), .S(n5842), .Z(n3891) );
  MUX2_X1 U5472 ( .A(n4991), .B(n6562), .S(n5842), .Z(n3890) );
  MUX2_X1 U5473 ( .A(n4992), .B(n6563), .S(n5842), .Z(n3889) );
  MUX2_X1 U5474 ( .A(n4993), .B(n6564), .S(n5842), .Z(n3888) );
  MUX2_X1 U5475 ( .A(n4994), .B(n6565), .S(n5842), .Z(n3887) );
  MUX2_X1 U5476 ( .A(n4995), .B(n6566), .S(n5842), .Z(n3886) );
  MUX2_X1 U5477 ( .A(n4996), .B(n6567), .S(n5842), .Z(n3885) );
  MUX2_X1 U5478 ( .A(n4997), .B(n6568), .S(n5842), .Z(n3884) );
  MUX2_X1 U5479 ( .A(n4998), .B(n6569), .S(n5842), .Z(n3883) );
  MUX2_X1 U5480 ( .A(n4999), .B(n6570), .S(n5842), .Z(n3882) );
  MUX2_X1 U5481 ( .A(n5000), .B(n6571), .S(n5842), .Z(n3881) );
  MUX2_X1 U5482 ( .A(n5001), .B(n6572), .S(n5842), .Z(n3880) );
  MUX2_X1 U5483 ( .A(n5002), .B(n6573), .S(n5842), .Z(n3879) );
  MUX2_X1 U5484 ( .A(n5003), .B(n6574), .S(n5842), .Z(n3878) );
  MUX2_X1 U5485 ( .A(n5004), .B(n6575), .S(n5842), .Z(n3877) );
  MUX2_X1 U5486 ( .A(n5005), .B(n6576), .S(n5842), .Z(n3876) );
  MUX2_X1 U5487 ( .A(n5006), .B(n6577), .S(n5842), .Z(n3875) );
  MUX2_X1 U5488 ( .A(n5007), .B(n6578), .S(n5842), .Z(n3874) );
  MUX2_X1 U5489 ( .A(n5008), .B(n6579), .S(n5842), .Z(n3873) );
  MUX2_X1 U5490 ( .A(n5009), .B(n6580), .S(n5842), .Z(n3872) );
  MUX2_X1 U5491 ( .A(n5010), .B(n6581), .S(n5842), .Z(n3871) );
  MUX2_X1 U5492 ( .A(n5011), .B(n6582), .S(n5842), .Z(n3870) );
  MUX2_X1 U5493 ( .A(n5012), .B(n6583), .S(n5842), .Z(n3869) );
  MUX2_X1 U5494 ( .A(n5013), .B(n6584), .S(n5842), .Z(n3868) );
  MUX2_X1 U5495 ( .A(n5014), .B(n6585), .S(n5842), .Z(n3867) );
  MUX2_X1 U5496 ( .A(n5015), .B(n6586), .S(n5842), .Z(n3866) );
  MUX2_X1 U5497 ( .A(n5016), .B(n6587), .S(n5842), .Z(n3865) );
  MUX2_X1 U5498 ( .A(n5017), .B(n6588), .S(n5842), .Z(n3864) );
  MUX2_X1 U5499 ( .A(n5018), .B(n6589), .S(n5842), .Z(n3863) );
  MUX2_X1 U5500 ( .A(n5019), .B(n6590), .S(n5842), .Z(n3862) );
  MUX2_X1 U5501 ( .A(n5020), .B(n6591), .S(n5842), .Z(n3861) );
  MUX2_X1 U5502 ( .A(n5021), .B(n6592), .S(n5842), .Z(n3860) );
  MUX2_X1 U5503 ( .A(n5022), .B(n6593), .S(n5842), .Z(n3859) );
  MUX2_X1 U5504 ( .A(n5023), .B(n6594), .S(n5842), .Z(n3858) );
  MUX2_X1 U5505 ( .A(n5024), .B(n6595), .S(n5842), .Z(n3857) );
  OAI211_X1 U5506 ( .C1(n6472), .C2(n6647), .A(n6650), .B(n6455), .ZN(n6649)
         );
  NAND3_X1 U5507 ( .A1(n6610), .A2(n6623), .A3(n6638), .ZN(n6650) );
  NOR2_X1 U5508 ( .A1(n6643), .A2(n6629), .ZN(n6610) );
  NAND2_X1 U5509 ( .A1(N208), .A2(n6651), .ZN(n6472) );
  MUX2_X1 U5510 ( .A(n6531), .B(n5236), .S(n6652), .Z(n3856) );
  MUX2_X1 U5511 ( .A(n6533), .B(n5237), .S(n6652), .Z(n3855) );
  MUX2_X1 U5512 ( .A(n6534), .B(n5238), .S(n6652), .Z(n3854) );
  MUX2_X1 U5513 ( .A(n6535), .B(n5239), .S(n6652), .Z(n3853) );
  MUX2_X1 U5514 ( .A(n6536), .B(n5240), .S(n6652), .Z(n3852) );
  MUX2_X1 U5515 ( .A(n6537), .B(n5241), .S(n6652), .Z(n3851) );
  MUX2_X1 U5516 ( .A(n6538), .B(n5242), .S(n6652), .Z(n3850) );
  MUX2_X1 U5517 ( .A(n6539), .B(n5243), .S(n6652), .Z(n3849) );
  MUX2_X1 U5518 ( .A(n6540), .B(n5244), .S(n6652), .Z(n3848) );
  MUX2_X1 U5519 ( .A(n6541), .B(n5245), .S(n6652), .Z(n3847) );
  MUX2_X1 U5520 ( .A(n6542), .B(n5246), .S(n6652), .Z(n3846) );
  MUX2_X1 U5521 ( .A(n6543), .B(n5247), .S(n6652), .Z(n3845) );
  MUX2_X1 U5522 ( .A(n6544), .B(n5248), .S(n6652), .Z(n3844) );
  MUX2_X1 U5523 ( .A(n6545), .B(n5249), .S(n6652), .Z(n3843) );
  MUX2_X1 U5524 ( .A(n6546), .B(n5250), .S(n6652), .Z(n3842) );
  MUX2_X1 U5525 ( .A(n6547), .B(n5251), .S(n6652), .Z(n3841) );
  MUX2_X1 U5526 ( .A(n6548), .B(n5252), .S(n6652), .Z(n3840) );
  MUX2_X1 U5527 ( .A(n6549), .B(n5253), .S(n6652), .Z(n3839) );
  MUX2_X1 U5528 ( .A(n6550), .B(n5254), .S(n6652), .Z(n3838) );
  MUX2_X1 U5529 ( .A(n6551), .B(n5255), .S(n6652), .Z(n3837) );
  MUX2_X1 U5530 ( .A(n6552), .B(n5256), .S(n6652), .Z(n3836) );
  MUX2_X1 U5531 ( .A(n6553), .B(n5257), .S(n6652), .Z(n3835) );
  MUX2_X1 U5532 ( .A(n6554), .B(n5258), .S(n6652), .Z(n3834) );
  MUX2_X1 U5533 ( .A(n6555), .B(n5259), .S(n6652), .Z(n3833) );
  MUX2_X1 U5534 ( .A(n6556), .B(n5260), .S(n6652), .Z(n3832) );
  MUX2_X1 U5535 ( .A(n6557), .B(n5261), .S(n6652), .Z(n3831) );
  MUX2_X1 U5536 ( .A(n6558), .B(n5262), .S(n6652), .Z(n3830) );
  MUX2_X1 U5537 ( .A(n6559), .B(n5263), .S(n6652), .Z(n3829) );
  MUX2_X1 U5538 ( .A(n6560), .B(n5264), .S(n6652), .Z(n3828) );
  MUX2_X1 U5539 ( .A(n6561), .B(n5265), .S(n6652), .Z(n3827) );
  MUX2_X1 U5540 ( .A(n6562), .B(n5266), .S(n6652), .Z(n3826) );
  MUX2_X1 U5541 ( .A(n6563), .B(n5267), .S(n6652), .Z(n3825) );
  MUX2_X1 U5542 ( .A(n6564), .B(n5268), .S(n6652), .Z(n3824) );
  MUX2_X1 U5543 ( .A(n6565), .B(n5269), .S(n6652), .Z(n3823) );
  MUX2_X1 U5544 ( .A(n6566), .B(n5270), .S(n6652), .Z(n3822) );
  MUX2_X1 U5545 ( .A(n6567), .B(n5271), .S(n6652), .Z(n3821) );
  MUX2_X1 U5546 ( .A(n6568), .B(n5272), .S(n6652), .Z(n3820) );
  MUX2_X1 U5547 ( .A(n6569), .B(n5273), .S(n6652), .Z(n3819) );
  MUX2_X1 U5548 ( .A(n6570), .B(n5274), .S(n6652), .Z(n3818) );
  MUX2_X1 U5549 ( .A(n6571), .B(n5275), .S(n6652), .Z(n3817) );
  MUX2_X1 U5550 ( .A(n6572), .B(n5276), .S(n6652), .Z(n3816) );
  MUX2_X1 U5551 ( .A(n6573), .B(n5277), .S(n6652), .Z(n3815) );
  MUX2_X1 U5552 ( .A(n6574), .B(n5278), .S(n6652), .Z(n3814) );
  MUX2_X1 U5553 ( .A(n6575), .B(n5279), .S(n6652), .Z(n3813) );
  MUX2_X1 U5554 ( .A(n6576), .B(n5280), .S(n6652), .Z(n3812) );
  MUX2_X1 U5555 ( .A(n6577), .B(n5281), .S(n6652), .Z(n3811) );
  MUX2_X1 U5556 ( .A(n6578), .B(n5282), .S(n6652), .Z(n3810) );
  MUX2_X1 U5557 ( .A(n6579), .B(n5283), .S(n6652), .Z(n3809) );
  MUX2_X1 U5558 ( .A(n6580), .B(n5284), .S(n6652), .Z(n3808) );
  MUX2_X1 U5559 ( .A(n6581), .B(n5285), .S(n6652), .Z(n3807) );
  MUX2_X1 U5560 ( .A(n6582), .B(n5286), .S(n6652), .Z(n3806) );
  MUX2_X1 U5561 ( .A(n6583), .B(n5287), .S(n6652), .Z(n3805) );
  MUX2_X1 U5562 ( .A(n6584), .B(n5288), .S(n6652), .Z(n3804) );
  MUX2_X1 U5563 ( .A(n6585), .B(n5289), .S(n6652), .Z(n3803) );
  MUX2_X1 U5564 ( .A(n6586), .B(n5290), .S(n6652), .Z(n3802) );
  MUX2_X1 U5565 ( .A(n6587), .B(n5291), .S(n6652), .Z(n3801) );
  MUX2_X1 U5566 ( .A(n6588), .B(n5292), .S(n6652), .Z(n3800) );
  MUX2_X1 U5567 ( .A(n6589), .B(n5293), .S(n6652), .Z(n3799) );
  MUX2_X1 U5568 ( .A(n6590), .B(n5294), .S(n6652), .Z(n3798) );
  MUX2_X1 U5569 ( .A(n6591), .B(n5295), .S(n6652), .Z(n3797) );
  MUX2_X1 U5570 ( .A(n6592), .B(n5296), .S(n6652), .Z(n3796) );
  MUX2_X1 U5571 ( .A(n6593), .B(n5297), .S(n6652), .Z(n3795) );
  MUX2_X1 U5572 ( .A(n6594), .B(n5298), .S(n6652), .Z(n3794) );
  MUX2_X1 U5573 ( .A(n6595), .B(n5299), .S(n6652), .Z(n3793) );
  INV_X1 U5574 ( .A(n6647), .ZN(n6653) );
  NAND2_X1 U5575 ( .A1(n6617), .A2(n6461), .ZN(n6647) );
  NOR2_X1 U5576 ( .A1(n6654), .A2(n5860), .ZN(n6617) );
  NOR2_X1 U5577 ( .A1(n6651), .A2(N208), .ZN(n6463) );
  AND2_X1 U5578 ( .A1(n6638), .A2(n6629), .ZN(n6635) );
  INV_X1 U5579 ( .A(n6655), .ZN(n6627) );
  MUX2_X1 U5580 ( .A(n6531), .B(n7988), .S(n6656), .Z(n3792) );
  INV_X1 U5581 ( .A(n6657), .ZN(n6531) );
  AOI22_X1 U5582 ( .A1(n5831), .A2(DATAIN[0]), .B1(n5834), .B2(BUSIN[0]), .ZN(
        n6657) );
  MUX2_X1 U5583 ( .A(n6533), .B(n7987), .S(n6656), .Z(n3791) );
  INV_X1 U5584 ( .A(n6658), .ZN(n6533) );
  AOI22_X1 U5585 ( .A1(n5831), .A2(DATAIN[1]), .B1(n5834), .B2(BUSIN[1]), .ZN(
        n6658) );
  MUX2_X1 U5586 ( .A(n6534), .B(n7986), .S(n6656), .Z(n3790) );
  INV_X1 U5587 ( .A(n6659), .ZN(n6534) );
  AOI22_X1 U5588 ( .A1(n5831), .A2(DATAIN[2]), .B1(n5834), .B2(BUSIN[2]), .ZN(
        n6659) );
  MUX2_X1 U5589 ( .A(n6535), .B(n7985), .S(n6656), .Z(n3789) );
  INV_X1 U5590 ( .A(n6660), .ZN(n6535) );
  AOI22_X1 U5591 ( .A1(n5831), .A2(DATAIN[3]), .B1(n5834), .B2(BUSIN[3]), .ZN(
        n6660) );
  MUX2_X1 U5592 ( .A(n6536), .B(n7984), .S(n6656), .Z(n3788) );
  INV_X1 U5593 ( .A(n6661), .ZN(n6536) );
  AOI22_X1 U5594 ( .A1(n5831), .A2(DATAIN[4]), .B1(n5834), .B2(BUSIN[4]), .ZN(
        n6661) );
  MUX2_X1 U5595 ( .A(n6537), .B(n7983), .S(n6656), .Z(n3787) );
  INV_X1 U5596 ( .A(n6662), .ZN(n6537) );
  AOI22_X1 U5597 ( .A1(n5831), .A2(DATAIN[5]), .B1(n5834), .B2(BUSIN[5]), .ZN(
        n6662) );
  MUX2_X1 U5598 ( .A(n6538), .B(n7982), .S(n6656), .Z(n3786) );
  INV_X1 U5599 ( .A(n6663), .ZN(n6538) );
  AOI22_X1 U5600 ( .A1(n5831), .A2(DATAIN[6]), .B1(n5834), .B2(BUSIN[6]), .ZN(
        n6663) );
  MUX2_X1 U5601 ( .A(n6539), .B(n7981), .S(n6656), .Z(n3785) );
  INV_X1 U5602 ( .A(n6664), .ZN(n6539) );
  AOI22_X1 U5603 ( .A1(n5831), .A2(DATAIN[7]), .B1(n5834), .B2(BUSIN[7]), .ZN(
        n6664) );
  MUX2_X1 U5604 ( .A(n6540), .B(n7980), .S(n6656), .Z(n3784) );
  INV_X1 U5605 ( .A(n6665), .ZN(n6540) );
  AOI22_X1 U5606 ( .A1(n5831), .A2(DATAIN[8]), .B1(n5834), .B2(BUSIN[8]), .ZN(
        n6665) );
  MUX2_X1 U5607 ( .A(n6541), .B(n7979), .S(n6656), .Z(n3783) );
  INV_X1 U5608 ( .A(n6666), .ZN(n6541) );
  AOI22_X1 U5609 ( .A1(n5831), .A2(DATAIN[9]), .B1(n5834), .B2(BUSIN[9]), .ZN(
        n6666) );
  MUX2_X1 U5610 ( .A(n6542), .B(n7978), .S(n6656), .Z(n3782) );
  INV_X1 U5611 ( .A(n6667), .ZN(n6542) );
  AOI22_X1 U5612 ( .A1(n5831), .A2(DATAIN[10]), .B1(n5834), .B2(BUSIN[10]), 
        .ZN(n6667) );
  MUX2_X1 U5613 ( .A(n6543), .B(n7977), .S(n6656), .Z(n3781) );
  INV_X1 U5614 ( .A(n6668), .ZN(n6543) );
  AOI22_X1 U5615 ( .A1(n5831), .A2(DATAIN[11]), .B1(n5834), .B2(BUSIN[11]), 
        .ZN(n6668) );
  MUX2_X1 U5616 ( .A(n6544), .B(n7976), .S(n6656), .Z(n3780) );
  INV_X1 U5617 ( .A(n6669), .ZN(n6544) );
  AOI22_X1 U5618 ( .A1(n5831), .A2(DATAIN[12]), .B1(n5834), .B2(BUSIN[12]), 
        .ZN(n6669) );
  MUX2_X1 U5619 ( .A(n6545), .B(n7975), .S(n6656), .Z(n3779) );
  INV_X1 U5620 ( .A(n6670), .ZN(n6545) );
  AOI22_X1 U5621 ( .A1(n5831), .A2(DATAIN[13]), .B1(n5834), .B2(BUSIN[13]), 
        .ZN(n6670) );
  MUX2_X1 U5622 ( .A(n6546), .B(n7974), .S(n6656), .Z(n3778) );
  INV_X1 U5623 ( .A(n6671), .ZN(n6546) );
  AOI22_X1 U5624 ( .A1(n5831), .A2(DATAIN[14]), .B1(n5834), .B2(BUSIN[14]), 
        .ZN(n6671) );
  MUX2_X1 U5625 ( .A(n6547), .B(n7973), .S(n6656), .Z(n3777) );
  INV_X1 U5626 ( .A(n6672), .ZN(n6547) );
  AOI22_X1 U5627 ( .A1(n5831), .A2(DATAIN[15]), .B1(n5834), .B2(BUSIN[15]), 
        .ZN(n6672) );
  MUX2_X1 U5628 ( .A(n6548), .B(n7972), .S(n6656), .Z(n3776) );
  INV_X1 U5629 ( .A(n6673), .ZN(n6548) );
  AOI22_X1 U5630 ( .A1(n5831), .A2(DATAIN[16]), .B1(n5834), .B2(BUSIN[16]), 
        .ZN(n6673) );
  MUX2_X1 U5631 ( .A(n6549), .B(n7971), .S(n6656), .Z(n3775) );
  INV_X1 U5632 ( .A(n6674), .ZN(n6549) );
  AOI22_X1 U5633 ( .A1(n5831), .A2(DATAIN[17]), .B1(n5834), .B2(BUSIN[17]), 
        .ZN(n6674) );
  MUX2_X1 U5634 ( .A(n6550), .B(n7970), .S(n6656), .Z(n3774) );
  INV_X1 U5635 ( .A(n6675), .ZN(n6550) );
  AOI22_X1 U5636 ( .A1(n5831), .A2(DATAIN[18]), .B1(n5834), .B2(BUSIN[18]), 
        .ZN(n6675) );
  MUX2_X1 U5637 ( .A(n6551), .B(n7969), .S(n6656), .Z(n3773) );
  INV_X1 U5638 ( .A(n6676), .ZN(n6551) );
  AOI22_X1 U5639 ( .A1(n5831), .A2(DATAIN[19]), .B1(n5834), .B2(BUSIN[19]), 
        .ZN(n6676) );
  MUX2_X1 U5640 ( .A(n6552), .B(n7968), .S(n6656), .Z(n3772) );
  INV_X1 U5641 ( .A(n6677), .ZN(n6552) );
  AOI22_X1 U5642 ( .A1(n5831), .A2(DATAIN[20]), .B1(n5834), .B2(BUSIN[20]), 
        .ZN(n6677) );
  MUX2_X1 U5643 ( .A(n6553), .B(n7967), .S(n6656), .Z(n3771) );
  INV_X1 U5644 ( .A(n6678), .ZN(n6553) );
  AOI22_X1 U5645 ( .A1(n5831), .A2(DATAIN[21]), .B1(n5834), .B2(BUSIN[21]), 
        .ZN(n6678) );
  MUX2_X1 U5646 ( .A(n6554), .B(n7966), .S(n6656), .Z(n3770) );
  INV_X1 U5647 ( .A(n6679), .ZN(n6554) );
  AOI22_X1 U5648 ( .A1(n5831), .A2(DATAIN[22]), .B1(n5834), .B2(BUSIN[22]), 
        .ZN(n6679) );
  MUX2_X1 U5649 ( .A(n6555), .B(n7965), .S(n6656), .Z(n3769) );
  INV_X1 U5650 ( .A(n6680), .ZN(n6555) );
  AOI22_X1 U5651 ( .A1(n5831), .A2(DATAIN[23]), .B1(n5834), .B2(BUSIN[23]), 
        .ZN(n6680) );
  MUX2_X1 U5652 ( .A(n6556), .B(n7964), .S(n6656), .Z(n3768) );
  INV_X1 U5653 ( .A(n6681), .ZN(n6556) );
  AOI22_X1 U5654 ( .A1(n5831), .A2(DATAIN[24]), .B1(n5834), .B2(BUSIN[24]), 
        .ZN(n6681) );
  MUX2_X1 U5655 ( .A(n6557), .B(n7963), .S(n6656), .Z(n3767) );
  INV_X1 U5656 ( .A(n6682), .ZN(n6557) );
  AOI22_X1 U5657 ( .A1(n5831), .A2(DATAIN[25]), .B1(n5834), .B2(BUSIN[25]), 
        .ZN(n6682) );
  MUX2_X1 U5658 ( .A(n6558), .B(n7962), .S(n6656), .Z(n3766) );
  INV_X1 U5659 ( .A(n6683), .ZN(n6558) );
  AOI22_X1 U5660 ( .A1(n5831), .A2(DATAIN[26]), .B1(n5834), .B2(BUSIN[26]), 
        .ZN(n6683) );
  MUX2_X1 U5661 ( .A(n6559), .B(n7961), .S(n6656), .Z(n3765) );
  INV_X1 U5662 ( .A(n6684), .ZN(n6559) );
  AOI22_X1 U5663 ( .A1(n5831), .A2(DATAIN[27]), .B1(n5834), .B2(BUSIN[27]), 
        .ZN(n6684) );
  MUX2_X1 U5664 ( .A(n6560), .B(n7960), .S(n6656), .Z(n3764) );
  INV_X1 U5665 ( .A(n6685), .ZN(n6560) );
  AOI22_X1 U5666 ( .A1(n5831), .A2(DATAIN[28]), .B1(n5834), .B2(BUSIN[28]), 
        .ZN(n6685) );
  MUX2_X1 U5667 ( .A(n6561), .B(n7959), .S(n6656), .Z(n3763) );
  INV_X1 U5668 ( .A(n6686), .ZN(n6561) );
  AOI22_X1 U5669 ( .A1(n5831), .A2(DATAIN[29]), .B1(n5834), .B2(BUSIN[29]), 
        .ZN(n6686) );
  MUX2_X1 U5670 ( .A(n6562), .B(n7958), .S(n6656), .Z(n3762) );
  INV_X1 U5671 ( .A(n6687), .ZN(n6562) );
  AOI22_X1 U5672 ( .A1(n5831), .A2(DATAIN[30]), .B1(n5834), .B2(BUSIN[30]), 
        .ZN(n6687) );
  MUX2_X1 U5673 ( .A(n6563), .B(n7957), .S(n6656), .Z(n3761) );
  INV_X1 U5674 ( .A(n6688), .ZN(n6563) );
  AOI22_X1 U5675 ( .A1(n5831), .A2(DATAIN[31]), .B1(n5834), .B2(BUSIN[31]), 
        .ZN(n6688) );
  MUX2_X1 U5676 ( .A(n6564), .B(n7956), .S(n6656), .Z(n3760) );
  INV_X1 U5677 ( .A(n6689), .ZN(n6564) );
  AOI22_X1 U5678 ( .A1(n5831), .A2(DATAIN[32]), .B1(n5834), .B2(BUSIN[32]), 
        .ZN(n6689) );
  MUX2_X1 U5679 ( .A(n6565), .B(n7955), .S(n6656), .Z(n3759) );
  INV_X1 U5680 ( .A(n6690), .ZN(n6565) );
  AOI22_X1 U5681 ( .A1(n5831), .A2(DATAIN[33]), .B1(n5834), .B2(BUSIN[33]), 
        .ZN(n6690) );
  MUX2_X1 U5682 ( .A(n6566), .B(n7954), .S(n6656), .Z(n3758) );
  INV_X1 U5683 ( .A(n6691), .ZN(n6566) );
  AOI22_X1 U5684 ( .A1(n5831), .A2(DATAIN[34]), .B1(n5834), .B2(BUSIN[34]), 
        .ZN(n6691) );
  MUX2_X1 U5685 ( .A(n6567), .B(n7953), .S(n6656), .Z(n3757) );
  INV_X1 U5686 ( .A(n6692), .ZN(n6567) );
  AOI22_X1 U5687 ( .A1(n5831), .A2(DATAIN[35]), .B1(n5834), .B2(BUSIN[35]), 
        .ZN(n6692) );
  MUX2_X1 U5688 ( .A(n6568), .B(n7952), .S(n6656), .Z(n3756) );
  INV_X1 U5689 ( .A(n6693), .ZN(n6568) );
  AOI22_X1 U5690 ( .A1(n5831), .A2(DATAIN[36]), .B1(n5834), .B2(BUSIN[36]), 
        .ZN(n6693) );
  MUX2_X1 U5691 ( .A(n6569), .B(n7951), .S(n6656), .Z(n3755) );
  INV_X1 U5692 ( .A(n6694), .ZN(n6569) );
  AOI22_X1 U5693 ( .A1(n5831), .A2(DATAIN[37]), .B1(n5834), .B2(BUSIN[37]), 
        .ZN(n6694) );
  MUX2_X1 U5694 ( .A(n6570), .B(n7950), .S(n6656), .Z(n3754) );
  INV_X1 U5695 ( .A(n6695), .ZN(n6570) );
  AOI22_X1 U5696 ( .A1(n5831), .A2(DATAIN[38]), .B1(n5834), .B2(BUSIN[38]), 
        .ZN(n6695) );
  MUX2_X1 U5697 ( .A(n6571), .B(n7949), .S(n6656), .Z(n3753) );
  INV_X1 U5698 ( .A(n6696), .ZN(n6571) );
  AOI22_X1 U5699 ( .A1(n5831), .A2(DATAIN[39]), .B1(n5834), .B2(BUSIN[39]), 
        .ZN(n6696) );
  MUX2_X1 U5700 ( .A(n6572), .B(n7948), .S(n6656), .Z(n3752) );
  INV_X1 U5701 ( .A(n6697), .ZN(n6572) );
  AOI22_X1 U5702 ( .A1(n5831), .A2(DATAIN[40]), .B1(n5834), .B2(BUSIN[40]), 
        .ZN(n6697) );
  MUX2_X1 U5703 ( .A(n6573), .B(n7947), .S(n6656), .Z(n3751) );
  INV_X1 U5704 ( .A(n6698), .ZN(n6573) );
  AOI22_X1 U5705 ( .A1(n5831), .A2(DATAIN[41]), .B1(n5834), .B2(BUSIN[41]), 
        .ZN(n6698) );
  MUX2_X1 U5706 ( .A(n6574), .B(n7946), .S(n6656), .Z(n3750) );
  INV_X1 U5707 ( .A(n6699), .ZN(n6574) );
  AOI22_X1 U5708 ( .A1(n5831), .A2(DATAIN[42]), .B1(n5834), .B2(BUSIN[42]), 
        .ZN(n6699) );
  MUX2_X1 U5709 ( .A(n6575), .B(n7945), .S(n6656), .Z(n3749) );
  INV_X1 U5710 ( .A(n6700), .ZN(n6575) );
  AOI22_X1 U5711 ( .A1(n5831), .A2(DATAIN[43]), .B1(n5834), .B2(BUSIN[43]), 
        .ZN(n6700) );
  MUX2_X1 U5712 ( .A(n6576), .B(n7944), .S(n6656), .Z(n3748) );
  INV_X1 U5713 ( .A(n6701), .ZN(n6576) );
  AOI22_X1 U5714 ( .A1(n5831), .A2(DATAIN[44]), .B1(n5834), .B2(BUSIN[44]), 
        .ZN(n6701) );
  MUX2_X1 U5715 ( .A(n6577), .B(n7943), .S(n6656), .Z(n3747) );
  INV_X1 U5716 ( .A(n6702), .ZN(n6577) );
  AOI22_X1 U5717 ( .A1(n5831), .A2(DATAIN[45]), .B1(n5834), .B2(BUSIN[45]), 
        .ZN(n6702) );
  MUX2_X1 U5718 ( .A(n6578), .B(n7942), .S(n6656), .Z(n3746) );
  INV_X1 U5719 ( .A(n6703), .ZN(n6578) );
  AOI22_X1 U5720 ( .A1(n5831), .A2(DATAIN[46]), .B1(n5834), .B2(BUSIN[46]), 
        .ZN(n6703) );
  MUX2_X1 U5721 ( .A(n6579), .B(n7941), .S(n6656), .Z(n3745) );
  INV_X1 U5722 ( .A(n6704), .ZN(n6579) );
  AOI22_X1 U5723 ( .A1(n5831), .A2(DATAIN[47]), .B1(n5834), .B2(BUSIN[47]), 
        .ZN(n6704) );
  MUX2_X1 U5724 ( .A(n6580), .B(n7940), .S(n6656), .Z(n3744) );
  INV_X1 U5725 ( .A(n6705), .ZN(n6580) );
  AOI22_X1 U5726 ( .A1(n5831), .A2(DATAIN[48]), .B1(n5834), .B2(BUSIN[48]), 
        .ZN(n6705) );
  MUX2_X1 U5727 ( .A(n6581), .B(n7939), .S(n6656), .Z(n3743) );
  INV_X1 U5728 ( .A(n6706), .ZN(n6581) );
  AOI22_X1 U5729 ( .A1(n5831), .A2(DATAIN[49]), .B1(n5834), .B2(BUSIN[49]), 
        .ZN(n6706) );
  MUX2_X1 U5730 ( .A(n6582), .B(n7938), .S(n6656), .Z(n3742) );
  INV_X1 U5731 ( .A(n6707), .ZN(n6582) );
  AOI22_X1 U5732 ( .A1(n5831), .A2(DATAIN[50]), .B1(n5834), .B2(BUSIN[50]), 
        .ZN(n6707) );
  MUX2_X1 U5733 ( .A(n6583), .B(n7937), .S(n6656), .Z(n3741) );
  INV_X1 U5734 ( .A(n6708), .ZN(n6583) );
  AOI22_X1 U5735 ( .A1(n5831), .A2(DATAIN[51]), .B1(n5834), .B2(BUSIN[51]), 
        .ZN(n6708) );
  MUX2_X1 U5736 ( .A(n6584), .B(n7936), .S(n6656), .Z(n3740) );
  INV_X1 U5737 ( .A(n6709), .ZN(n6584) );
  AOI22_X1 U5738 ( .A1(n5831), .A2(DATAIN[52]), .B1(n5834), .B2(BUSIN[52]), 
        .ZN(n6709) );
  MUX2_X1 U5739 ( .A(n6585), .B(n7935), .S(n6656), .Z(n3739) );
  INV_X1 U5740 ( .A(n6710), .ZN(n6585) );
  AOI22_X1 U5741 ( .A1(n5831), .A2(DATAIN[53]), .B1(n5834), .B2(BUSIN[53]), 
        .ZN(n6710) );
  MUX2_X1 U5742 ( .A(n6586), .B(n7934), .S(n6656), .Z(n3738) );
  INV_X1 U5743 ( .A(n6711), .ZN(n6586) );
  AOI22_X1 U5744 ( .A1(n5831), .A2(DATAIN[54]), .B1(n5834), .B2(BUSIN[54]), 
        .ZN(n6711) );
  MUX2_X1 U5745 ( .A(n6587), .B(n7933), .S(n6656), .Z(n3737) );
  INV_X1 U5746 ( .A(n6712), .ZN(n6587) );
  AOI22_X1 U5747 ( .A1(n5831), .A2(DATAIN[55]), .B1(n5834), .B2(BUSIN[55]), 
        .ZN(n6712) );
  MUX2_X1 U5748 ( .A(n6588), .B(n7932), .S(n6656), .Z(n3736) );
  INV_X1 U5749 ( .A(n6713), .ZN(n6588) );
  AOI22_X1 U5750 ( .A1(n5831), .A2(DATAIN[56]), .B1(n5834), .B2(BUSIN[56]), 
        .ZN(n6713) );
  MUX2_X1 U5751 ( .A(n6589), .B(n7931), .S(n6656), .Z(n3735) );
  INV_X1 U5752 ( .A(n6714), .ZN(n6589) );
  AOI22_X1 U5753 ( .A1(n5831), .A2(DATAIN[57]), .B1(n5834), .B2(BUSIN[57]), 
        .ZN(n6714) );
  MUX2_X1 U5754 ( .A(n6590), .B(n7930), .S(n6656), .Z(n3734) );
  INV_X1 U5755 ( .A(n6715), .ZN(n6590) );
  AOI22_X1 U5756 ( .A1(n5831), .A2(DATAIN[58]), .B1(n5834), .B2(BUSIN[58]), 
        .ZN(n6715) );
  MUX2_X1 U5757 ( .A(n6591), .B(n7929), .S(n6656), .Z(n3733) );
  INV_X1 U5758 ( .A(n6716), .ZN(n6591) );
  AOI22_X1 U5759 ( .A1(n5831), .A2(DATAIN[59]), .B1(n5834), .B2(BUSIN[59]), 
        .ZN(n6716) );
  MUX2_X1 U5760 ( .A(n6592), .B(n7928), .S(n6656), .Z(n3732) );
  INV_X1 U5761 ( .A(n6717), .ZN(n6592) );
  AOI22_X1 U5762 ( .A1(n5831), .A2(DATAIN[60]), .B1(n5834), .B2(BUSIN[60]), 
        .ZN(n6717) );
  MUX2_X1 U5763 ( .A(n6593), .B(n7927), .S(n6656), .Z(n3731) );
  INV_X1 U5764 ( .A(n6718), .ZN(n6593) );
  AOI22_X1 U5765 ( .A1(n5831), .A2(DATAIN[61]), .B1(n5834), .B2(BUSIN[61]), 
        .ZN(n6718) );
  MUX2_X1 U5766 ( .A(n6594), .B(n7926), .S(n6656), .Z(n3730) );
  INV_X1 U5767 ( .A(n6719), .ZN(n6594) );
  AOI22_X1 U5768 ( .A1(n5831), .A2(DATAIN[62]), .B1(n5834), .B2(BUSIN[62]), 
        .ZN(n6719) );
  MUX2_X1 U5769 ( .A(n6595), .B(n7925), .S(n6656), .Z(n3729) );
  NOR2_X1 U5770 ( .A1(n6631), .A2(n6598), .ZN(n6638) );
  NOR2_X1 U5771 ( .A1(n6655), .A2(n6629), .ZN(n6600) );
  NAND2_X1 U5772 ( .A1(n6623), .A2(n6643), .ZN(n6655) );
  NOR2_X1 U5773 ( .A1(n6720), .A2(n6644), .ZN(n6623) );
  NOR2_X1 U5774 ( .A1(N210), .A2(N209), .ZN(n6461) );
  NOR2_X1 U5775 ( .A1(n5855), .A2(N208), .ZN(n6467) );
  INV_X1 U5776 ( .A(n6721), .ZN(n6595) );
  AOI22_X1 U5777 ( .A1(n5831), .A2(DATAIN[63]), .B1(n5834), .B2(BUSIN[63]), 
        .ZN(n6721) );
  NAND4_X1 U5778 ( .A1(n6722), .A2(n6723), .A3(n6724), .A4(n6725), .ZN(n3728)
         );
  AOI221_X1 U5779 ( .B1(n6726), .B2(n5236), .C1(n6727), .C2(n4961), .A(n6728), 
        .ZN(n6725) );
  OAI222_X1 U5780 ( .A1(n1121), .A2(n5821), .B1(n1057), .B2(n5828), .C1(n1185), 
        .C2(n5817), .ZN(n6728) );
  AOI221_X1 U5781 ( .B1(n6729), .B2(n5301), .C1(n6730), .C2(n5090), .A(n6731), 
        .ZN(n6724) );
  OAI222_X1 U5782 ( .A1(n609), .A2(n6732), .B1(n545), .B2(n5829), .C1(n801), 
        .C2(n6733), .ZN(n6731) );
  AOI221_X1 U5783 ( .B1(n6734), .B2(n8180), .C1(n6735), .C2(n8116), .A(n6736), 
        .ZN(n6723) );
  OAI222_X1 U5784 ( .A1(n5026), .A2(n6737), .B1(n993), .B2(n5822), .C1(n5429), 
        .C2(n5818), .ZN(n6736) );
  AOI221_X1 U5785 ( .B1(n5832), .B2(DATAIN[0]), .C1(n6738), .C2(OUT1[0]), .A(
        n6739), .ZN(n6722) );
  OAI22_X1 U5786 ( .A1(n4831), .A2(n5826), .B1(n5365), .B2(n6740), .ZN(n6739)
         );
  NAND4_X1 U5787 ( .A1(n6741), .A2(n6742), .A3(n6743), .A4(n6744), .ZN(n3727)
         );
  AOI221_X1 U5788 ( .B1(n6726), .B2(n5237), .C1(n6727), .C2(n4962), .A(n6745), 
        .ZN(n6744) );
  OAI222_X1 U5789 ( .A1(n1120), .A2(n5821), .B1(n1056), .B2(n5828), .C1(n1184), 
        .C2(n5817), .ZN(n6745) );
  AOI221_X1 U5790 ( .B1(n6729), .B2(n5302), .C1(n6730), .C2(n5091), .A(n6746), 
        .ZN(n6743) );
  OAI222_X1 U5791 ( .A1(n608), .A2(n6732), .B1(n544), .B2(n5829), .C1(n800), 
        .C2(n6733), .ZN(n6746) );
  AOI221_X1 U5792 ( .B1(n6734), .B2(n8179), .C1(n6735), .C2(n8115), .A(n6747), 
        .ZN(n6742) );
  OAI222_X1 U5793 ( .A1(n5027), .A2(n6737), .B1(n992), .B2(n5822), .C1(n5430), 
        .C2(n5818), .ZN(n6747) );
  AOI221_X1 U5794 ( .B1(n5832), .B2(DATAIN[1]), .C1(n6738), .C2(OUT1[1]), .A(
        n6748), .ZN(n6741) );
  OAI22_X1 U5795 ( .A1(n4832), .A2(n5826), .B1(n5366), .B2(n6740), .ZN(n6748)
         );
  NAND4_X1 U5796 ( .A1(n6749), .A2(n6750), .A3(n6751), .A4(n6752), .ZN(n3726)
         );
  AOI221_X1 U5797 ( .B1(n6726), .B2(n5238), .C1(n6727), .C2(n4963), .A(n6753), 
        .ZN(n6752) );
  OAI222_X1 U5798 ( .A1(n1119), .A2(n5821), .B1(n1055), .B2(n5828), .C1(n1183), 
        .C2(n5817), .ZN(n6753) );
  AOI221_X1 U5799 ( .B1(n6729), .B2(n5303), .C1(n6730), .C2(n5092), .A(n6754), 
        .ZN(n6751) );
  OAI222_X1 U5800 ( .A1(n607), .A2(n6732), .B1(n543), .B2(n5829), .C1(n799), 
        .C2(n6733), .ZN(n6754) );
  AOI221_X1 U5801 ( .B1(n6734), .B2(n8178), .C1(n6735), .C2(n8114), .A(n6755), 
        .ZN(n6750) );
  OAI222_X1 U5802 ( .A1(n5028), .A2(n6737), .B1(n991), .B2(n5822), .C1(n5431), 
        .C2(n5818), .ZN(n6755) );
  AOI221_X1 U5803 ( .B1(n5832), .B2(DATAIN[2]), .C1(n6738), .C2(OUT1[2]), .A(
        n6756), .ZN(n6749) );
  OAI22_X1 U5804 ( .A1(n4833), .A2(n5826), .B1(n5367), .B2(n6740), .ZN(n6756)
         );
  NAND4_X1 U5805 ( .A1(n6757), .A2(n6758), .A3(n6759), .A4(n6760), .ZN(n3725)
         );
  AOI221_X1 U5806 ( .B1(n6726), .B2(n5239), .C1(n6727), .C2(n4964), .A(n6761), 
        .ZN(n6760) );
  OAI222_X1 U5807 ( .A1(n1118), .A2(n5821), .B1(n1054), .B2(n5828), .C1(n1182), 
        .C2(n5817), .ZN(n6761) );
  AOI221_X1 U5808 ( .B1(n6729), .B2(n5304), .C1(n6730), .C2(n5093), .A(n6762), 
        .ZN(n6759) );
  OAI222_X1 U5809 ( .A1(n606), .A2(n6732), .B1(n542), .B2(n5829), .C1(n798), 
        .C2(n6733), .ZN(n6762) );
  AOI221_X1 U5810 ( .B1(n6734), .B2(n8177), .C1(n6735), .C2(n8113), .A(n6763), 
        .ZN(n6758) );
  OAI222_X1 U5811 ( .A1(n5029), .A2(n6737), .B1(n990), .B2(n5822), .C1(n5432), 
        .C2(n5818), .ZN(n6763) );
  AOI221_X1 U5812 ( .B1(n5832), .B2(DATAIN[3]), .C1(n6738), .C2(OUT1[3]), .A(
        n6764), .ZN(n6757) );
  OAI22_X1 U5813 ( .A1(n4834), .A2(n5826), .B1(n5368), .B2(n6740), .ZN(n6764)
         );
  NAND4_X1 U5814 ( .A1(n6765), .A2(n6766), .A3(n6767), .A4(n6768), .ZN(n3724)
         );
  AOI221_X1 U5815 ( .B1(n6726), .B2(n5240), .C1(n6727), .C2(n4965), .A(n6769), 
        .ZN(n6768) );
  OAI222_X1 U5816 ( .A1(n1117), .A2(n5821), .B1(n1053), .B2(n5828), .C1(n1181), 
        .C2(n5817), .ZN(n6769) );
  AOI221_X1 U5817 ( .B1(n6729), .B2(n5305), .C1(n6730), .C2(n5094), .A(n6770), 
        .ZN(n6767) );
  OAI222_X1 U5818 ( .A1(n605), .A2(n6732), .B1(n541), .B2(n5829), .C1(n797), 
        .C2(n6733), .ZN(n6770) );
  AOI221_X1 U5819 ( .B1(n6734), .B2(n8176), .C1(n6735), .C2(n8112), .A(n6771), 
        .ZN(n6766) );
  OAI222_X1 U5820 ( .A1(n5030), .A2(n6737), .B1(n989), .B2(n5822), .C1(n5433), 
        .C2(n5818), .ZN(n6771) );
  AOI221_X1 U5821 ( .B1(n5832), .B2(DATAIN[4]), .C1(n6738), .C2(OUT1[4]), .A(
        n6772), .ZN(n6765) );
  OAI22_X1 U5822 ( .A1(n4835), .A2(n5826), .B1(n5369), .B2(n6740), .ZN(n6772)
         );
  NAND4_X1 U5823 ( .A1(n6773), .A2(n6774), .A3(n6775), .A4(n6776), .ZN(n3723)
         );
  AOI221_X1 U5824 ( .B1(n6726), .B2(n5241), .C1(n6727), .C2(n4966), .A(n6777), 
        .ZN(n6776) );
  OAI222_X1 U5825 ( .A1(n1116), .A2(n5821), .B1(n1052), .B2(n5828), .C1(n1180), 
        .C2(n5817), .ZN(n6777) );
  AOI221_X1 U5826 ( .B1(n6729), .B2(n5306), .C1(n6730), .C2(n5095), .A(n6778), 
        .ZN(n6775) );
  OAI222_X1 U5827 ( .A1(n604), .A2(n6732), .B1(n540), .B2(n5829), .C1(n796), 
        .C2(n6733), .ZN(n6778) );
  AOI221_X1 U5828 ( .B1(n6734), .B2(n8175), .C1(n6735), .C2(n8111), .A(n6779), 
        .ZN(n6774) );
  OAI222_X1 U5829 ( .A1(n5031), .A2(n6737), .B1(n988), .B2(n5822), .C1(n5434), 
        .C2(n5818), .ZN(n6779) );
  AOI221_X1 U5830 ( .B1(n5832), .B2(DATAIN[5]), .C1(n6738), .C2(OUT1[5]), .A(
        n6780), .ZN(n6773) );
  OAI22_X1 U5831 ( .A1(n4836), .A2(n5826), .B1(n5370), .B2(n6740), .ZN(n6780)
         );
  NAND4_X1 U5832 ( .A1(n6781), .A2(n6782), .A3(n6783), .A4(n6784), .ZN(n3722)
         );
  AOI221_X1 U5833 ( .B1(n6726), .B2(n5242), .C1(n6727), .C2(n4967), .A(n6785), 
        .ZN(n6784) );
  OAI222_X1 U5834 ( .A1(n1115), .A2(n5821), .B1(n1051), .B2(n5828), .C1(n1179), 
        .C2(n5817), .ZN(n6785) );
  AOI221_X1 U5835 ( .B1(n6729), .B2(n5307), .C1(n6730), .C2(n5096), .A(n6786), 
        .ZN(n6783) );
  OAI222_X1 U5836 ( .A1(n603), .A2(n6732), .B1(n539), .B2(n5829), .C1(n795), 
        .C2(n6733), .ZN(n6786) );
  AOI221_X1 U5837 ( .B1(n6734), .B2(n8174), .C1(n6735), .C2(n8110), .A(n6787), 
        .ZN(n6782) );
  OAI222_X1 U5838 ( .A1(n5032), .A2(n6737), .B1(n987), .B2(n5822), .C1(n5435), 
        .C2(n5818), .ZN(n6787) );
  AOI221_X1 U5839 ( .B1(n5832), .B2(DATAIN[6]), .C1(n6738), .C2(OUT1[6]), .A(
        n6788), .ZN(n6781) );
  OAI22_X1 U5840 ( .A1(n4837), .A2(n5826), .B1(n5371), .B2(n6740), .ZN(n6788)
         );
  NAND4_X1 U5841 ( .A1(n6789), .A2(n6790), .A3(n6791), .A4(n6792), .ZN(n3721)
         );
  AOI221_X1 U5842 ( .B1(n6726), .B2(n5243), .C1(n6727), .C2(n4968), .A(n6793), 
        .ZN(n6792) );
  OAI222_X1 U5843 ( .A1(n1114), .A2(n5821), .B1(n1050), .B2(n5828), .C1(n1178), 
        .C2(n5817), .ZN(n6793) );
  AOI221_X1 U5844 ( .B1(n6729), .B2(n5308), .C1(n6730), .C2(n5097), .A(n6794), 
        .ZN(n6791) );
  OAI222_X1 U5845 ( .A1(n602), .A2(n6732), .B1(n538), .B2(n5829), .C1(n794), 
        .C2(n6733), .ZN(n6794) );
  AOI221_X1 U5846 ( .B1(n6734), .B2(n8173), .C1(n6735), .C2(n8109), .A(n6795), 
        .ZN(n6790) );
  OAI222_X1 U5847 ( .A1(n5033), .A2(n6737), .B1(n986), .B2(n5822), .C1(n5436), 
        .C2(n5818), .ZN(n6795) );
  AOI221_X1 U5848 ( .B1(n5832), .B2(DATAIN[7]), .C1(n6738), .C2(OUT1[7]), .A(
        n6796), .ZN(n6789) );
  OAI22_X1 U5849 ( .A1(n4838), .A2(n5826), .B1(n5372), .B2(n6740), .ZN(n6796)
         );
  NAND4_X1 U5850 ( .A1(n6797), .A2(n6798), .A3(n6799), .A4(n6800), .ZN(n3720)
         );
  AOI221_X1 U5851 ( .B1(n6726), .B2(n5244), .C1(n6727), .C2(n4969), .A(n6801), 
        .ZN(n6800) );
  OAI222_X1 U5852 ( .A1(n1113), .A2(n5821), .B1(n1049), .B2(n5828), .C1(n1177), 
        .C2(n5817), .ZN(n6801) );
  AOI221_X1 U5853 ( .B1(n6729), .B2(n5309), .C1(n6730), .C2(n5098), .A(n6802), 
        .ZN(n6799) );
  OAI222_X1 U5854 ( .A1(n601), .A2(n6732), .B1(n537), .B2(n5829), .C1(n793), 
        .C2(n6733), .ZN(n6802) );
  AOI221_X1 U5855 ( .B1(n6734), .B2(n8172), .C1(n6735), .C2(n8108), .A(n6803), 
        .ZN(n6798) );
  OAI222_X1 U5856 ( .A1(n5034), .A2(n6737), .B1(n985), .B2(n5822), .C1(n5437), 
        .C2(n5818), .ZN(n6803) );
  AOI221_X1 U5857 ( .B1(n5832), .B2(DATAIN[8]), .C1(n6738), .C2(OUT1[8]), .A(
        n6804), .ZN(n6797) );
  OAI22_X1 U5858 ( .A1(n4839), .A2(n5826), .B1(n5373), .B2(n6740), .ZN(n6804)
         );
  NAND4_X1 U5859 ( .A1(n6805), .A2(n6806), .A3(n6807), .A4(n6808), .ZN(n3719)
         );
  AOI221_X1 U5860 ( .B1(n6726), .B2(n5245), .C1(n6727), .C2(n4970), .A(n6809), 
        .ZN(n6808) );
  OAI222_X1 U5861 ( .A1(n1112), .A2(n5821), .B1(n1048), .B2(n5828), .C1(n1176), 
        .C2(n5817), .ZN(n6809) );
  AOI221_X1 U5862 ( .B1(n6729), .B2(n5310), .C1(n6730), .C2(n5099), .A(n6810), 
        .ZN(n6807) );
  OAI222_X1 U5863 ( .A1(n600), .A2(n6732), .B1(n536), .B2(n5829), .C1(n792), 
        .C2(n6733), .ZN(n6810) );
  AOI221_X1 U5864 ( .B1(n6734), .B2(n8171), .C1(n6735), .C2(n8107), .A(n6811), 
        .ZN(n6806) );
  OAI222_X1 U5865 ( .A1(n5035), .A2(n6737), .B1(n984), .B2(n5822), .C1(n5438), 
        .C2(n5818), .ZN(n6811) );
  AOI221_X1 U5866 ( .B1(n5832), .B2(DATAIN[9]), .C1(n6738), .C2(OUT1[9]), .A(
        n6812), .ZN(n6805) );
  OAI22_X1 U5867 ( .A1(n4840), .A2(n5826), .B1(n5374), .B2(n6740), .ZN(n6812)
         );
  NAND4_X1 U5868 ( .A1(n6813), .A2(n6814), .A3(n6815), .A4(n6816), .ZN(n3718)
         );
  AOI221_X1 U5869 ( .B1(n6726), .B2(n5246), .C1(n6727), .C2(n4971), .A(n6817), 
        .ZN(n6816) );
  OAI222_X1 U5870 ( .A1(n1111), .A2(n5821), .B1(n1047), .B2(n5828), .C1(n1175), 
        .C2(n5817), .ZN(n6817) );
  AOI221_X1 U5871 ( .B1(n6729), .B2(n5311), .C1(n6730), .C2(n5100), .A(n6818), 
        .ZN(n6815) );
  OAI222_X1 U5872 ( .A1(n599), .A2(n6732), .B1(n535), .B2(n5829), .C1(n791), 
        .C2(n6733), .ZN(n6818) );
  AOI221_X1 U5873 ( .B1(n6734), .B2(n8170), .C1(n6735), .C2(n8106), .A(n6819), 
        .ZN(n6814) );
  OAI222_X1 U5874 ( .A1(n5036), .A2(n6737), .B1(n983), .B2(n5822), .C1(n5439), 
        .C2(n5818), .ZN(n6819) );
  AOI221_X1 U5875 ( .B1(n5832), .B2(DATAIN[10]), .C1(n6738), .C2(OUT1[10]), 
        .A(n6820), .ZN(n6813) );
  OAI22_X1 U5876 ( .A1(n4841), .A2(n5826), .B1(n5375), .B2(n6740), .ZN(n6820)
         );
  NAND4_X1 U5877 ( .A1(n6821), .A2(n6822), .A3(n6823), .A4(n6824), .ZN(n3717)
         );
  AOI221_X1 U5878 ( .B1(n6726), .B2(n5247), .C1(n6727), .C2(n4972), .A(n6825), 
        .ZN(n6824) );
  OAI222_X1 U5879 ( .A1(n1110), .A2(n5821), .B1(n1046), .B2(n5828), .C1(n1174), 
        .C2(n5817), .ZN(n6825) );
  AOI221_X1 U5880 ( .B1(n6729), .B2(n5312), .C1(n6730), .C2(n5101), .A(n6826), 
        .ZN(n6823) );
  OAI222_X1 U5881 ( .A1(n598), .A2(n6732), .B1(n534), .B2(n5829), .C1(n790), 
        .C2(n6733), .ZN(n6826) );
  AOI221_X1 U5882 ( .B1(n6734), .B2(n8169), .C1(n6735), .C2(n8105), .A(n6827), 
        .ZN(n6822) );
  OAI222_X1 U5883 ( .A1(n5037), .A2(n6737), .B1(n982), .B2(n5822), .C1(n5440), 
        .C2(n5818), .ZN(n6827) );
  AOI221_X1 U5884 ( .B1(n5832), .B2(DATAIN[11]), .C1(n6738), .C2(OUT1[11]), 
        .A(n6828), .ZN(n6821) );
  OAI22_X1 U5885 ( .A1(n4842), .A2(n5826), .B1(n5376), .B2(n6740), .ZN(n6828)
         );
  NAND4_X1 U5886 ( .A1(n6829), .A2(n6830), .A3(n6831), .A4(n6832), .ZN(n3716)
         );
  AOI221_X1 U5887 ( .B1(n6726), .B2(n5248), .C1(n6727), .C2(n4973), .A(n6833), 
        .ZN(n6832) );
  OAI222_X1 U5888 ( .A1(n1109), .A2(n5821), .B1(n1045), .B2(n5828), .C1(n1173), 
        .C2(n5817), .ZN(n6833) );
  AOI221_X1 U5889 ( .B1(n6729), .B2(n5313), .C1(n6730), .C2(n5102), .A(n6834), 
        .ZN(n6831) );
  OAI222_X1 U5890 ( .A1(n597), .A2(n6732), .B1(n533), .B2(n5829), .C1(n789), 
        .C2(n6733), .ZN(n6834) );
  AOI221_X1 U5891 ( .B1(n6734), .B2(n8168), .C1(n6735), .C2(n8104), .A(n6835), 
        .ZN(n6830) );
  OAI222_X1 U5892 ( .A1(n5038), .A2(n6737), .B1(n981), .B2(n5822), .C1(n5441), 
        .C2(n5818), .ZN(n6835) );
  AOI221_X1 U5893 ( .B1(n5832), .B2(DATAIN[12]), .C1(n6738), .C2(OUT1[12]), 
        .A(n6836), .ZN(n6829) );
  OAI22_X1 U5894 ( .A1(n4843), .A2(n5826), .B1(n5377), .B2(n6740), .ZN(n6836)
         );
  NAND4_X1 U5895 ( .A1(n6837), .A2(n6838), .A3(n6839), .A4(n6840), .ZN(n3715)
         );
  AOI221_X1 U5896 ( .B1(n6726), .B2(n5249), .C1(n6727), .C2(n4974), .A(n6841), 
        .ZN(n6840) );
  OAI222_X1 U5897 ( .A1(n1108), .A2(n5821), .B1(n1044), .B2(n5828), .C1(n1172), 
        .C2(n5817), .ZN(n6841) );
  AOI221_X1 U5898 ( .B1(n6729), .B2(n5314), .C1(n6730), .C2(n5103), .A(n6842), 
        .ZN(n6839) );
  OAI222_X1 U5899 ( .A1(n596), .A2(n6732), .B1(n532), .B2(n5829), .C1(n788), 
        .C2(n6733), .ZN(n6842) );
  AOI221_X1 U5900 ( .B1(n6734), .B2(n8167), .C1(n6735), .C2(n8103), .A(n6843), 
        .ZN(n6838) );
  OAI222_X1 U5901 ( .A1(n5039), .A2(n6737), .B1(n980), .B2(n5822), .C1(n5442), 
        .C2(n5818), .ZN(n6843) );
  AOI221_X1 U5902 ( .B1(n5832), .B2(DATAIN[13]), .C1(n6738), .C2(OUT1[13]), 
        .A(n6844), .ZN(n6837) );
  OAI22_X1 U5903 ( .A1(n4844), .A2(n5826), .B1(n5378), .B2(n6740), .ZN(n6844)
         );
  NAND4_X1 U5904 ( .A1(n6845), .A2(n6846), .A3(n6847), .A4(n6848), .ZN(n3714)
         );
  AOI221_X1 U5905 ( .B1(n6726), .B2(n5250), .C1(n6727), .C2(n4975), .A(n6849), 
        .ZN(n6848) );
  OAI222_X1 U5906 ( .A1(n1107), .A2(n5821), .B1(n1043), .B2(n5828), .C1(n1171), 
        .C2(n5817), .ZN(n6849) );
  AOI221_X1 U5907 ( .B1(n6729), .B2(n5315), .C1(n6730), .C2(n5104), .A(n6850), 
        .ZN(n6847) );
  OAI222_X1 U5908 ( .A1(n595), .A2(n6732), .B1(n531), .B2(n5829), .C1(n787), 
        .C2(n6733), .ZN(n6850) );
  AOI221_X1 U5909 ( .B1(n6734), .B2(n8166), .C1(n6735), .C2(n8102), .A(n6851), 
        .ZN(n6846) );
  OAI222_X1 U5910 ( .A1(n5040), .A2(n6737), .B1(n979), .B2(n5822), .C1(n5443), 
        .C2(n5818), .ZN(n6851) );
  AOI221_X1 U5911 ( .B1(n5832), .B2(DATAIN[14]), .C1(n6738), .C2(OUT1[14]), 
        .A(n6852), .ZN(n6845) );
  OAI22_X1 U5912 ( .A1(n4845), .A2(n5826), .B1(n5379), .B2(n6740), .ZN(n6852)
         );
  NAND4_X1 U5913 ( .A1(n6853), .A2(n6854), .A3(n6855), .A4(n6856), .ZN(n3713)
         );
  AOI221_X1 U5914 ( .B1(n6726), .B2(n5251), .C1(n6727), .C2(n4976), .A(n6857), 
        .ZN(n6856) );
  OAI222_X1 U5915 ( .A1(n1106), .A2(n5821), .B1(n1042), .B2(n5828), .C1(n1170), 
        .C2(n5817), .ZN(n6857) );
  AOI221_X1 U5916 ( .B1(n6729), .B2(n5316), .C1(n6730), .C2(n5105), .A(n6858), 
        .ZN(n6855) );
  OAI222_X1 U5917 ( .A1(n594), .A2(n6732), .B1(n530), .B2(n5829), .C1(n786), 
        .C2(n6733), .ZN(n6858) );
  AOI221_X1 U5918 ( .B1(n6734), .B2(n8165), .C1(n6735), .C2(n8101), .A(n6859), 
        .ZN(n6854) );
  OAI222_X1 U5919 ( .A1(n5041), .A2(n6737), .B1(n978), .B2(n5822), .C1(n5444), 
        .C2(n5818), .ZN(n6859) );
  AOI221_X1 U5920 ( .B1(n5832), .B2(DATAIN[15]), .C1(n6738), .C2(OUT1[15]), 
        .A(n6860), .ZN(n6853) );
  OAI22_X1 U5921 ( .A1(n4846), .A2(n5826), .B1(n5380), .B2(n6740), .ZN(n6860)
         );
  NAND4_X1 U5922 ( .A1(n6861), .A2(n6862), .A3(n6863), .A4(n6864), .ZN(n3712)
         );
  AOI221_X1 U5923 ( .B1(n6726), .B2(n5252), .C1(n6727), .C2(n4977), .A(n6865), 
        .ZN(n6864) );
  OAI222_X1 U5924 ( .A1(n1105), .A2(n5821), .B1(n1041), .B2(n5828), .C1(n1169), 
        .C2(n5817), .ZN(n6865) );
  AOI221_X1 U5925 ( .B1(n6729), .B2(n5317), .C1(n6730), .C2(n5106), .A(n6866), 
        .ZN(n6863) );
  OAI222_X1 U5926 ( .A1(n593), .A2(n6732), .B1(n529), .B2(n5829), .C1(n785), 
        .C2(n6733), .ZN(n6866) );
  AOI221_X1 U5927 ( .B1(n6734), .B2(n8164), .C1(n6735), .C2(n8100), .A(n6867), 
        .ZN(n6862) );
  OAI222_X1 U5928 ( .A1(n5042), .A2(n6737), .B1(n977), .B2(n5822), .C1(n5445), 
        .C2(n5818), .ZN(n6867) );
  AOI221_X1 U5929 ( .B1(n5832), .B2(DATAIN[16]), .C1(n6738), .C2(OUT1[16]), 
        .A(n6868), .ZN(n6861) );
  OAI22_X1 U5930 ( .A1(n4847), .A2(n5826), .B1(n5381), .B2(n6740), .ZN(n6868)
         );
  NAND4_X1 U5931 ( .A1(n6869), .A2(n6870), .A3(n6871), .A4(n6872), .ZN(n3711)
         );
  AOI221_X1 U5932 ( .B1(n6726), .B2(n5253), .C1(n6727), .C2(n4978), .A(n6873), 
        .ZN(n6872) );
  OAI222_X1 U5933 ( .A1(n1104), .A2(n5821), .B1(n1040), .B2(n5828), .C1(n1168), 
        .C2(n5817), .ZN(n6873) );
  AOI221_X1 U5934 ( .B1(n6729), .B2(n5318), .C1(n6730), .C2(n5107), .A(n6874), 
        .ZN(n6871) );
  OAI222_X1 U5935 ( .A1(n592), .A2(n6732), .B1(n528), .B2(n5829), .C1(n784), 
        .C2(n6733), .ZN(n6874) );
  AOI221_X1 U5936 ( .B1(n6734), .B2(n8163), .C1(n6735), .C2(n8099), .A(n6875), 
        .ZN(n6870) );
  OAI222_X1 U5937 ( .A1(n5043), .A2(n6737), .B1(n976), .B2(n5822), .C1(n5446), 
        .C2(n5818), .ZN(n6875) );
  AOI221_X1 U5938 ( .B1(n5832), .B2(DATAIN[17]), .C1(n6738), .C2(OUT1[17]), 
        .A(n6876), .ZN(n6869) );
  OAI22_X1 U5939 ( .A1(n4848), .A2(n5826), .B1(n5382), .B2(n6740), .ZN(n6876)
         );
  NAND4_X1 U5940 ( .A1(n6877), .A2(n6878), .A3(n6879), .A4(n6880), .ZN(n3710)
         );
  AOI221_X1 U5941 ( .B1(n6726), .B2(n5254), .C1(n6727), .C2(n4979), .A(n6881), 
        .ZN(n6880) );
  OAI222_X1 U5942 ( .A1(n1103), .A2(n5821), .B1(n1039), .B2(n5828), .C1(n1167), 
        .C2(n5817), .ZN(n6881) );
  AOI221_X1 U5943 ( .B1(n6729), .B2(n5319), .C1(n6730), .C2(n5108), .A(n6882), 
        .ZN(n6879) );
  OAI222_X1 U5944 ( .A1(n591), .A2(n6732), .B1(n527), .B2(n5829), .C1(n783), 
        .C2(n6733), .ZN(n6882) );
  AOI221_X1 U5945 ( .B1(n6734), .B2(n8162), .C1(n6735), .C2(n8098), .A(n6883), 
        .ZN(n6878) );
  OAI222_X1 U5946 ( .A1(n5044), .A2(n6737), .B1(n975), .B2(n5822), .C1(n5447), 
        .C2(n5818), .ZN(n6883) );
  AOI221_X1 U5947 ( .B1(n5832), .B2(DATAIN[18]), .C1(n6738), .C2(OUT1[18]), 
        .A(n6884), .ZN(n6877) );
  OAI22_X1 U5948 ( .A1(n4849), .A2(n5826), .B1(n5383), .B2(n6740), .ZN(n6884)
         );
  NAND4_X1 U5949 ( .A1(n6885), .A2(n6886), .A3(n6887), .A4(n6888), .ZN(n3709)
         );
  AOI221_X1 U5950 ( .B1(n6726), .B2(n5255), .C1(n6727), .C2(n4980), .A(n6889), 
        .ZN(n6888) );
  OAI222_X1 U5951 ( .A1(n1102), .A2(n5821), .B1(n1038), .B2(n5828), .C1(n1166), 
        .C2(n5817), .ZN(n6889) );
  AOI221_X1 U5952 ( .B1(n6729), .B2(n5320), .C1(n6730), .C2(n5109), .A(n6890), 
        .ZN(n6887) );
  OAI222_X1 U5953 ( .A1(n590), .A2(n6732), .B1(n526), .B2(n5829), .C1(n782), 
        .C2(n6733), .ZN(n6890) );
  AOI221_X1 U5954 ( .B1(n6734), .B2(n8161), .C1(n6735), .C2(n8097), .A(n6891), 
        .ZN(n6886) );
  OAI222_X1 U5955 ( .A1(n5045), .A2(n6737), .B1(n974), .B2(n5822), .C1(n5448), 
        .C2(n5818), .ZN(n6891) );
  AOI221_X1 U5956 ( .B1(n5832), .B2(DATAIN[19]), .C1(n6738), .C2(OUT1[19]), 
        .A(n6892), .ZN(n6885) );
  OAI22_X1 U5957 ( .A1(n4850), .A2(n5826), .B1(n5384), .B2(n6740), .ZN(n6892)
         );
  NAND4_X1 U5958 ( .A1(n6893), .A2(n6894), .A3(n6895), .A4(n6896), .ZN(n3708)
         );
  AOI221_X1 U5959 ( .B1(n6726), .B2(n5256), .C1(n6727), .C2(n4981), .A(n6897), 
        .ZN(n6896) );
  OAI222_X1 U5960 ( .A1(n1101), .A2(n5821), .B1(n1037), .B2(n5828), .C1(n1165), 
        .C2(n5817), .ZN(n6897) );
  AOI221_X1 U5961 ( .B1(n6729), .B2(n5321), .C1(n6730), .C2(n5110), .A(n6898), 
        .ZN(n6895) );
  OAI222_X1 U5962 ( .A1(n589), .A2(n6732), .B1(n525), .B2(n5829), .C1(n781), 
        .C2(n6733), .ZN(n6898) );
  AOI221_X1 U5963 ( .B1(n6734), .B2(n8160), .C1(n6735), .C2(n8096), .A(n6899), 
        .ZN(n6894) );
  OAI222_X1 U5964 ( .A1(n5046), .A2(n6737), .B1(n973), .B2(n5822), .C1(n5449), 
        .C2(n5818), .ZN(n6899) );
  AOI221_X1 U5965 ( .B1(n5832), .B2(DATAIN[20]), .C1(n6738), .C2(OUT1[20]), 
        .A(n6900), .ZN(n6893) );
  OAI22_X1 U5966 ( .A1(n4851), .A2(n5826), .B1(n5385), .B2(n6740), .ZN(n6900)
         );
  NAND4_X1 U5967 ( .A1(n6901), .A2(n6902), .A3(n6903), .A4(n6904), .ZN(n3707)
         );
  AOI221_X1 U5968 ( .B1(n6726), .B2(n5257), .C1(n6727), .C2(n4982), .A(n6905), 
        .ZN(n6904) );
  OAI222_X1 U5969 ( .A1(n1100), .A2(n5821), .B1(n1036), .B2(n5828), .C1(n1164), 
        .C2(n5817), .ZN(n6905) );
  AOI221_X1 U5970 ( .B1(n6729), .B2(n5322), .C1(n6730), .C2(n5111), .A(n6906), 
        .ZN(n6903) );
  OAI222_X1 U5971 ( .A1(n588), .A2(n6732), .B1(n524), .B2(n5829), .C1(n780), 
        .C2(n6733), .ZN(n6906) );
  AOI221_X1 U5972 ( .B1(n6734), .B2(n8159), .C1(n6735), .C2(n8095), .A(n6907), 
        .ZN(n6902) );
  OAI222_X1 U5973 ( .A1(n5047), .A2(n6737), .B1(n972), .B2(n5822), .C1(n5450), 
        .C2(n5818), .ZN(n6907) );
  AOI221_X1 U5974 ( .B1(n5832), .B2(DATAIN[21]), .C1(n6738), .C2(OUT1[21]), 
        .A(n6908), .ZN(n6901) );
  OAI22_X1 U5975 ( .A1(n4852), .A2(n5826), .B1(n5386), .B2(n6740), .ZN(n6908)
         );
  NAND4_X1 U5976 ( .A1(n6909), .A2(n6910), .A3(n6911), .A4(n6912), .ZN(n3706)
         );
  AOI221_X1 U5977 ( .B1(n6726), .B2(n5258), .C1(n6727), .C2(n4983), .A(n6913), 
        .ZN(n6912) );
  OAI222_X1 U5978 ( .A1(n1099), .A2(n5821), .B1(n1035), .B2(n5828), .C1(n1163), 
        .C2(n5817), .ZN(n6913) );
  AOI221_X1 U5979 ( .B1(n6729), .B2(n5323), .C1(n6730), .C2(n5112), .A(n6914), 
        .ZN(n6911) );
  OAI222_X1 U5980 ( .A1(n587), .A2(n6732), .B1(n523), .B2(n5829), .C1(n779), 
        .C2(n6733), .ZN(n6914) );
  AOI221_X1 U5981 ( .B1(n6734), .B2(n8158), .C1(n6735), .C2(n8094), .A(n6915), 
        .ZN(n6910) );
  OAI222_X1 U5982 ( .A1(n5048), .A2(n6737), .B1(n971), .B2(n5822), .C1(n5451), 
        .C2(n5818), .ZN(n6915) );
  AOI221_X1 U5983 ( .B1(n5832), .B2(DATAIN[22]), .C1(n6738), .C2(OUT1[22]), 
        .A(n6916), .ZN(n6909) );
  OAI22_X1 U5984 ( .A1(n4853), .A2(n5826), .B1(n5387), .B2(n6740), .ZN(n6916)
         );
  NAND4_X1 U5985 ( .A1(n6917), .A2(n6918), .A3(n6919), .A4(n6920), .ZN(n3705)
         );
  AOI221_X1 U5986 ( .B1(n6726), .B2(n5259), .C1(n6727), .C2(n4984), .A(n6921), 
        .ZN(n6920) );
  OAI222_X1 U5987 ( .A1(n1098), .A2(n5821), .B1(n1034), .B2(n5828), .C1(n1162), 
        .C2(n5817), .ZN(n6921) );
  AOI221_X1 U5988 ( .B1(n6729), .B2(n5324), .C1(n6730), .C2(n5113), .A(n6922), 
        .ZN(n6919) );
  OAI222_X1 U5989 ( .A1(n586), .A2(n6732), .B1(n522), .B2(n5829), .C1(n778), 
        .C2(n6733), .ZN(n6922) );
  AOI221_X1 U5990 ( .B1(n6734), .B2(n8157), .C1(n6735), .C2(n8093), .A(n6923), 
        .ZN(n6918) );
  OAI222_X1 U5991 ( .A1(n5049), .A2(n6737), .B1(n970), .B2(n5822), .C1(n5452), 
        .C2(n5818), .ZN(n6923) );
  AOI221_X1 U5992 ( .B1(n5832), .B2(DATAIN[23]), .C1(n6738), .C2(OUT1[23]), 
        .A(n6924), .ZN(n6917) );
  OAI22_X1 U5993 ( .A1(n4854), .A2(n5826), .B1(n5388), .B2(n6740), .ZN(n6924)
         );
  NAND4_X1 U5994 ( .A1(n6925), .A2(n6926), .A3(n6927), .A4(n6928), .ZN(n3704)
         );
  AOI221_X1 U5995 ( .B1(n6726), .B2(n5260), .C1(n6727), .C2(n4985), .A(n6929), 
        .ZN(n6928) );
  OAI222_X1 U5996 ( .A1(n1097), .A2(n5821), .B1(n1033), .B2(n5828), .C1(n1161), 
        .C2(n5817), .ZN(n6929) );
  AOI221_X1 U5997 ( .B1(n6729), .B2(n5325), .C1(n6730), .C2(n5114), .A(n6930), 
        .ZN(n6927) );
  OAI222_X1 U5998 ( .A1(n585), .A2(n6732), .B1(n521), .B2(n5829), .C1(n777), 
        .C2(n6733), .ZN(n6930) );
  AOI221_X1 U5999 ( .B1(n6734), .B2(n8156), .C1(n6735), .C2(n8092), .A(n6931), 
        .ZN(n6926) );
  OAI222_X1 U6000 ( .A1(n5050), .A2(n6737), .B1(n969), .B2(n5822), .C1(n5453), 
        .C2(n5818), .ZN(n6931) );
  AOI221_X1 U6001 ( .B1(n5832), .B2(DATAIN[24]), .C1(n6738), .C2(OUT1[24]), 
        .A(n6932), .ZN(n6925) );
  OAI22_X1 U6002 ( .A1(n4855), .A2(n5826), .B1(n5389), .B2(n6740), .ZN(n6932)
         );
  NAND4_X1 U6003 ( .A1(n6933), .A2(n6934), .A3(n6935), .A4(n6936), .ZN(n3703)
         );
  AOI221_X1 U6004 ( .B1(n6726), .B2(n5261), .C1(n6727), .C2(n4986), .A(n6937), 
        .ZN(n6936) );
  OAI222_X1 U6005 ( .A1(n1096), .A2(n5821), .B1(n1032), .B2(n5828), .C1(n1160), 
        .C2(n5817), .ZN(n6937) );
  AOI221_X1 U6006 ( .B1(n6729), .B2(n5326), .C1(n6730), .C2(n5115), .A(n6938), 
        .ZN(n6935) );
  OAI222_X1 U6007 ( .A1(n584), .A2(n6732), .B1(n520), .B2(n5829), .C1(n776), 
        .C2(n6733), .ZN(n6938) );
  AOI221_X1 U6008 ( .B1(n6734), .B2(n8155), .C1(n6735), .C2(n8091), .A(n6939), 
        .ZN(n6934) );
  OAI222_X1 U6009 ( .A1(n5051), .A2(n6737), .B1(n968), .B2(n5822), .C1(n5454), 
        .C2(n5818), .ZN(n6939) );
  AOI221_X1 U6010 ( .B1(n5832), .B2(DATAIN[25]), .C1(n6738), .C2(OUT1[25]), 
        .A(n6940), .ZN(n6933) );
  OAI22_X1 U6011 ( .A1(n4856), .A2(n5826), .B1(n5390), .B2(n6740), .ZN(n6940)
         );
  NAND4_X1 U6012 ( .A1(n6941), .A2(n6942), .A3(n6943), .A4(n6944), .ZN(n3702)
         );
  AOI221_X1 U6013 ( .B1(n6726), .B2(n5262), .C1(n6727), .C2(n4987), .A(n6945), 
        .ZN(n6944) );
  OAI222_X1 U6014 ( .A1(n1095), .A2(n5821), .B1(n1031), .B2(n5828), .C1(n1159), 
        .C2(n5817), .ZN(n6945) );
  AOI221_X1 U6015 ( .B1(n6729), .B2(n5327), .C1(n6730), .C2(n5116), .A(n6946), 
        .ZN(n6943) );
  OAI222_X1 U6016 ( .A1(n583), .A2(n6732), .B1(n519), .B2(n5829), .C1(n775), 
        .C2(n6733), .ZN(n6946) );
  AOI221_X1 U6017 ( .B1(n6734), .B2(n8154), .C1(n6735), .C2(n8090), .A(n6947), 
        .ZN(n6942) );
  OAI222_X1 U6018 ( .A1(n5052), .A2(n6737), .B1(n967), .B2(n5822), .C1(n5455), 
        .C2(n5818), .ZN(n6947) );
  AOI221_X1 U6019 ( .B1(n5832), .B2(DATAIN[26]), .C1(n6738), .C2(OUT1[26]), 
        .A(n6948), .ZN(n6941) );
  OAI22_X1 U6020 ( .A1(n4857), .A2(n5826), .B1(n5391), .B2(n6740), .ZN(n6948)
         );
  NAND4_X1 U6021 ( .A1(n6949), .A2(n6950), .A3(n6951), .A4(n6952), .ZN(n3701)
         );
  AOI221_X1 U6022 ( .B1(n6726), .B2(n5263), .C1(n6727), .C2(n4988), .A(n6953), 
        .ZN(n6952) );
  OAI222_X1 U6023 ( .A1(n1094), .A2(n5821), .B1(n1030), .B2(n5828), .C1(n1158), 
        .C2(n5817), .ZN(n6953) );
  AOI221_X1 U6024 ( .B1(n6729), .B2(n5328), .C1(n6730), .C2(n5117), .A(n6954), 
        .ZN(n6951) );
  OAI222_X1 U6025 ( .A1(n582), .A2(n6732), .B1(n518), .B2(n5829), .C1(n774), 
        .C2(n6733), .ZN(n6954) );
  AOI221_X1 U6026 ( .B1(n6734), .B2(n8153), .C1(n6735), .C2(n8089), .A(n6955), 
        .ZN(n6950) );
  OAI222_X1 U6027 ( .A1(n5053), .A2(n6737), .B1(n966), .B2(n5822), .C1(n5456), 
        .C2(n5818), .ZN(n6955) );
  AOI221_X1 U6028 ( .B1(n5832), .B2(DATAIN[27]), .C1(n6738), .C2(OUT1[27]), 
        .A(n6956), .ZN(n6949) );
  OAI22_X1 U6029 ( .A1(n4858), .A2(n5826), .B1(n5392), .B2(n6740), .ZN(n6956)
         );
  NAND4_X1 U6030 ( .A1(n6957), .A2(n6958), .A3(n6959), .A4(n6960), .ZN(n3700)
         );
  AOI221_X1 U6031 ( .B1(n6726), .B2(n5264), .C1(n6727), .C2(n4989), .A(n6961), 
        .ZN(n6960) );
  OAI222_X1 U6032 ( .A1(n1093), .A2(n5821), .B1(n1029), .B2(n5828), .C1(n1157), 
        .C2(n5817), .ZN(n6961) );
  AOI221_X1 U6033 ( .B1(n6729), .B2(n5329), .C1(n6730), .C2(n5118), .A(n6962), 
        .ZN(n6959) );
  OAI222_X1 U6034 ( .A1(n581), .A2(n6732), .B1(n517), .B2(n5829), .C1(n773), 
        .C2(n6733), .ZN(n6962) );
  AOI221_X1 U6035 ( .B1(n6734), .B2(n8152), .C1(n6735), .C2(n8088), .A(n6963), 
        .ZN(n6958) );
  OAI222_X1 U6036 ( .A1(n5054), .A2(n6737), .B1(n965), .B2(n5822), .C1(n5457), 
        .C2(n5818), .ZN(n6963) );
  AOI221_X1 U6037 ( .B1(n5832), .B2(DATAIN[28]), .C1(n6738), .C2(OUT1[28]), 
        .A(n6964), .ZN(n6957) );
  OAI22_X1 U6038 ( .A1(n4859), .A2(n5826), .B1(n5393), .B2(n6740), .ZN(n6964)
         );
  NAND4_X1 U6039 ( .A1(n6965), .A2(n6966), .A3(n6967), .A4(n6968), .ZN(n3699)
         );
  AOI221_X1 U6040 ( .B1(n6726), .B2(n5265), .C1(n6727), .C2(n4990), .A(n6969), 
        .ZN(n6968) );
  OAI222_X1 U6041 ( .A1(n1092), .A2(n5821), .B1(n1028), .B2(n5828), .C1(n1156), 
        .C2(n5817), .ZN(n6969) );
  AOI221_X1 U6042 ( .B1(n6729), .B2(n5330), .C1(n6730), .C2(n5119), .A(n6970), 
        .ZN(n6967) );
  OAI222_X1 U6043 ( .A1(n580), .A2(n6732), .B1(n516), .B2(n5829), .C1(n772), 
        .C2(n6733), .ZN(n6970) );
  AOI221_X1 U6044 ( .B1(n6734), .B2(n8151), .C1(n6735), .C2(n8087), .A(n6971), 
        .ZN(n6966) );
  OAI222_X1 U6045 ( .A1(n5055), .A2(n6737), .B1(n964), .B2(n5822), .C1(n5458), 
        .C2(n5818), .ZN(n6971) );
  AOI221_X1 U6046 ( .B1(n5832), .B2(DATAIN[29]), .C1(n6738), .C2(OUT1[29]), 
        .A(n6972), .ZN(n6965) );
  OAI22_X1 U6047 ( .A1(n4860), .A2(n5826), .B1(n5394), .B2(n6740), .ZN(n6972)
         );
  NAND4_X1 U6048 ( .A1(n6973), .A2(n6974), .A3(n6975), .A4(n6976), .ZN(n3698)
         );
  AOI221_X1 U6049 ( .B1(n6726), .B2(n5266), .C1(n6727), .C2(n4991), .A(n6977), 
        .ZN(n6976) );
  OAI222_X1 U6050 ( .A1(n1091), .A2(n5821), .B1(n1027), .B2(n5828), .C1(n1155), 
        .C2(n5817), .ZN(n6977) );
  AOI221_X1 U6051 ( .B1(n6729), .B2(n5331), .C1(n6730), .C2(n5120), .A(n6978), 
        .ZN(n6975) );
  OAI222_X1 U6052 ( .A1(n579), .A2(n6732), .B1(n515), .B2(n5829), .C1(n771), 
        .C2(n6733), .ZN(n6978) );
  AOI221_X1 U6053 ( .B1(n6734), .B2(n8150), .C1(n6735), .C2(n8086), .A(n6979), 
        .ZN(n6974) );
  OAI222_X1 U6054 ( .A1(n5056), .A2(n6737), .B1(n963), .B2(n5822), .C1(n5459), 
        .C2(n5818), .ZN(n6979) );
  AOI221_X1 U6055 ( .B1(n5832), .B2(DATAIN[30]), .C1(n6738), .C2(OUT1[30]), 
        .A(n6980), .ZN(n6973) );
  OAI22_X1 U6056 ( .A1(n4861), .A2(n5826), .B1(n5395), .B2(n6740), .ZN(n6980)
         );
  NAND4_X1 U6057 ( .A1(n6981), .A2(n6982), .A3(n6983), .A4(n6984), .ZN(n3697)
         );
  AOI221_X1 U6058 ( .B1(n6726), .B2(n5267), .C1(n6727), .C2(n4992), .A(n6985), 
        .ZN(n6984) );
  OAI222_X1 U6059 ( .A1(n1090), .A2(n5821), .B1(n1026), .B2(n5828), .C1(n1154), 
        .C2(n5817), .ZN(n6985) );
  AOI221_X1 U6060 ( .B1(n6729), .B2(n5332), .C1(n6730), .C2(n5121), .A(n6986), 
        .ZN(n6983) );
  OAI222_X1 U6061 ( .A1(n578), .A2(n6732), .B1(n514), .B2(n5829), .C1(n770), 
        .C2(n6733), .ZN(n6986) );
  AOI221_X1 U6062 ( .B1(n6734), .B2(n8149), .C1(n6735), .C2(n8085), .A(n6987), 
        .ZN(n6982) );
  OAI222_X1 U6063 ( .A1(n5057), .A2(n6737), .B1(n962), .B2(n5822), .C1(n5460), 
        .C2(n5818), .ZN(n6987) );
  AOI221_X1 U6064 ( .B1(n5832), .B2(DATAIN[31]), .C1(n6738), .C2(OUT1[31]), 
        .A(n6988), .ZN(n6981) );
  OAI22_X1 U6065 ( .A1(n4862), .A2(n5826), .B1(n5396), .B2(n6740), .ZN(n6988)
         );
  NAND4_X1 U6066 ( .A1(n6989), .A2(n6990), .A3(n6991), .A4(n6992), .ZN(n3696)
         );
  AOI221_X1 U6067 ( .B1(n6726), .B2(n5268), .C1(n6727), .C2(n4993), .A(n6993), 
        .ZN(n6992) );
  OAI222_X1 U6068 ( .A1(n1089), .A2(n5821), .B1(n1025), .B2(n5828), .C1(n1153), 
        .C2(n5817), .ZN(n6993) );
  AOI221_X1 U6069 ( .B1(n6729), .B2(n5333), .C1(n6730), .C2(n5122), .A(n6994), 
        .ZN(n6991) );
  OAI222_X1 U6070 ( .A1(n577), .A2(n6732), .B1(n513), .B2(n5829), .C1(n769), 
        .C2(n6733), .ZN(n6994) );
  AOI221_X1 U6071 ( .B1(n6734), .B2(n8148), .C1(n6735), .C2(n8084), .A(n6995), 
        .ZN(n6990) );
  OAI222_X1 U6072 ( .A1(n5058), .A2(n6737), .B1(n961), .B2(n5822), .C1(n5461), 
        .C2(n5818), .ZN(n6995) );
  AOI221_X1 U6073 ( .B1(n5832), .B2(DATAIN[32]), .C1(n6738), .C2(OUT1[32]), 
        .A(n6996), .ZN(n6989) );
  OAI22_X1 U6074 ( .A1(n4863), .A2(n5826), .B1(n5397), .B2(n6740), .ZN(n6996)
         );
  NAND4_X1 U6075 ( .A1(n6997), .A2(n6998), .A3(n6999), .A4(n7000), .ZN(n3695)
         );
  AOI221_X1 U6076 ( .B1(n6726), .B2(n5269), .C1(n6727), .C2(n4994), .A(n7001), 
        .ZN(n7000) );
  OAI222_X1 U6077 ( .A1(n1088), .A2(n5821), .B1(n1024), .B2(n5828), .C1(n1152), 
        .C2(n5817), .ZN(n7001) );
  AOI221_X1 U6078 ( .B1(n6729), .B2(n5334), .C1(n6730), .C2(n5123), .A(n7002), 
        .ZN(n6999) );
  OAI222_X1 U6079 ( .A1(n576), .A2(n6732), .B1(n512), .B2(n5829), .C1(n768), 
        .C2(n6733), .ZN(n7002) );
  AOI221_X1 U6080 ( .B1(n6734), .B2(n8147), .C1(n6735), .C2(n8083), .A(n7003), 
        .ZN(n6998) );
  OAI222_X1 U6081 ( .A1(n5059), .A2(n6737), .B1(n960), .B2(n5822), .C1(n5462), 
        .C2(n5818), .ZN(n7003) );
  AOI221_X1 U6082 ( .B1(n5832), .B2(DATAIN[33]), .C1(n6738), .C2(OUT1[33]), 
        .A(n7004), .ZN(n6997) );
  OAI22_X1 U6083 ( .A1(n4864), .A2(n5826), .B1(n5398), .B2(n6740), .ZN(n7004)
         );
  NAND4_X1 U6084 ( .A1(n7005), .A2(n7006), .A3(n7007), .A4(n7008), .ZN(n3694)
         );
  AOI221_X1 U6085 ( .B1(n6726), .B2(n5270), .C1(n6727), .C2(n4995), .A(n7009), 
        .ZN(n7008) );
  OAI222_X1 U6086 ( .A1(n1087), .A2(n5821), .B1(n1023), .B2(n5828), .C1(n1151), 
        .C2(n5817), .ZN(n7009) );
  AOI221_X1 U6087 ( .B1(n6729), .B2(n5335), .C1(n6730), .C2(n5124), .A(n7010), 
        .ZN(n7007) );
  OAI222_X1 U6088 ( .A1(n575), .A2(n6732), .B1(n511), .B2(n5829), .C1(n767), 
        .C2(n6733), .ZN(n7010) );
  AOI221_X1 U6089 ( .B1(n6734), .B2(n8146), .C1(n6735), .C2(n8082), .A(n7011), 
        .ZN(n7006) );
  OAI222_X1 U6090 ( .A1(n5060), .A2(n6737), .B1(n959), .B2(n5822), .C1(n5463), 
        .C2(n5818), .ZN(n7011) );
  AOI221_X1 U6091 ( .B1(n5832), .B2(DATAIN[34]), .C1(n6738), .C2(OUT1[34]), 
        .A(n7012), .ZN(n7005) );
  OAI22_X1 U6092 ( .A1(n4865), .A2(n5826), .B1(n5399), .B2(n6740), .ZN(n7012)
         );
  NAND4_X1 U6093 ( .A1(n7013), .A2(n7014), .A3(n7015), .A4(n7016), .ZN(n3693)
         );
  AOI221_X1 U6094 ( .B1(n6726), .B2(n5271), .C1(n6727), .C2(n4996), .A(n7017), 
        .ZN(n7016) );
  OAI222_X1 U6095 ( .A1(n1086), .A2(n5821), .B1(n1022), .B2(n5828), .C1(n1150), 
        .C2(n5817), .ZN(n7017) );
  AOI221_X1 U6096 ( .B1(n6729), .B2(n5336), .C1(n6730), .C2(n5125), .A(n7018), 
        .ZN(n7015) );
  OAI222_X1 U6097 ( .A1(n574), .A2(n6732), .B1(n510), .B2(n5829), .C1(n766), 
        .C2(n6733), .ZN(n7018) );
  AOI221_X1 U6098 ( .B1(n6734), .B2(n8145), .C1(n6735), .C2(n8081), .A(n7019), 
        .ZN(n7014) );
  OAI222_X1 U6099 ( .A1(n5061), .A2(n6737), .B1(n958), .B2(n5822), .C1(n5464), 
        .C2(n5818), .ZN(n7019) );
  AOI221_X1 U6100 ( .B1(n5832), .B2(DATAIN[35]), .C1(n6738), .C2(OUT1[35]), 
        .A(n7020), .ZN(n7013) );
  OAI22_X1 U6101 ( .A1(n4866), .A2(n5826), .B1(n5400), .B2(n6740), .ZN(n7020)
         );
  NAND4_X1 U6102 ( .A1(n7021), .A2(n7022), .A3(n7023), .A4(n7024), .ZN(n3692)
         );
  AOI221_X1 U6103 ( .B1(n6726), .B2(n5272), .C1(n6727), .C2(n4997), .A(n7025), 
        .ZN(n7024) );
  OAI222_X1 U6104 ( .A1(n1085), .A2(n5821), .B1(n1021), .B2(n5828), .C1(n1149), 
        .C2(n5817), .ZN(n7025) );
  AOI221_X1 U6105 ( .B1(n6729), .B2(n5337), .C1(n6730), .C2(n5126), .A(n7026), 
        .ZN(n7023) );
  OAI222_X1 U6106 ( .A1(n573), .A2(n6732), .B1(n509), .B2(n5829), .C1(n765), 
        .C2(n6733), .ZN(n7026) );
  AOI221_X1 U6107 ( .B1(n6734), .B2(n8144), .C1(n6735), .C2(n8080), .A(n7027), 
        .ZN(n7022) );
  OAI222_X1 U6108 ( .A1(n5062), .A2(n6737), .B1(n957), .B2(n5822), .C1(n5465), 
        .C2(n5818), .ZN(n7027) );
  AOI221_X1 U6109 ( .B1(n5832), .B2(DATAIN[36]), .C1(n6738), .C2(OUT1[36]), 
        .A(n7028), .ZN(n7021) );
  OAI22_X1 U6110 ( .A1(n4867), .A2(n5826), .B1(n5401), .B2(n6740), .ZN(n7028)
         );
  NAND4_X1 U6111 ( .A1(n7029), .A2(n7030), .A3(n7031), .A4(n7032), .ZN(n3691)
         );
  AOI221_X1 U6112 ( .B1(n6726), .B2(n5273), .C1(n6727), .C2(n4998), .A(n7033), 
        .ZN(n7032) );
  OAI222_X1 U6113 ( .A1(n1084), .A2(n5821), .B1(n1020), .B2(n5828), .C1(n1148), 
        .C2(n5817), .ZN(n7033) );
  AOI221_X1 U6114 ( .B1(n6729), .B2(n5338), .C1(n6730), .C2(n5127), .A(n7034), 
        .ZN(n7031) );
  OAI222_X1 U6115 ( .A1(n572), .A2(n6732), .B1(n508), .B2(n5829), .C1(n764), 
        .C2(n6733), .ZN(n7034) );
  AOI221_X1 U6116 ( .B1(n6734), .B2(n8143), .C1(n6735), .C2(n8079), .A(n7035), 
        .ZN(n7030) );
  OAI222_X1 U6117 ( .A1(n5063), .A2(n6737), .B1(n956), .B2(n5822), .C1(n5466), 
        .C2(n5818), .ZN(n7035) );
  AOI221_X1 U6118 ( .B1(n5832), .B2(DATAIN[37]), .C1(n6738), .C2(OUT1[37]), 
        .A(n7036), .ZN(n7029) );
  OAI22_X1 U6119 ( .A1(n4868), .A2(n5826), .B1(n5402), .B2(n6740), .ZN(n7036)
         );
  NAND4_X1 U6120 ( .A1(n7037), .A2(n7038), .A3(n7039), .A4(n7040), .ZN(n3690)
         );
  AOI221_X1 U6121 ( .B1(n6726), .B2(n5274), .C1(n6727), .C2(n4999), .A(n7041), 
        .ZN(n7040) );
  OAI222_X1 U6122 ( .A1(n1083), .A2(n5821), .B1(n1019), .B2(n5828), .C1(n1147), 
        .C2(n5817), .ZN(n7041) );
  AOI221_X1 U6123 ( .B1(n6729), .B2(n5339), .C1(n6730), .C2(n5128), .A(n7042), 
        .ZN(n7039) );
  OAI222_X1 U6124 ( .A1(n571), .A2(n6732), .B1(n507), .B2(n5829), .C1(n763), 
        .C2(n6733), .ZN(n7042) );
  AOI221_X1 U6125 ( .B1(n6734), .B2(n8142), .C1(n6735), .C2(n8078), .A(n7043), 
        .ZN(n7038) );
  OAI222_X1 U6126 ( .A1(n5064), .A2(n6737), .B1(n955), .B2(n5822), .C1(n5467), 
        .C2(n5818), .ZN(n7043) );
  AOI221_X1 U6127 ( .B1(n5832), .B2(DATAIN[38]), .C1(n6738), .C2(OUT1[38]), 
        .A(n7044), .ZN(n7037) );
  OAI22_X1 U6128 ( .A1(n4869), .A2(n5826), .B1(n5403), .B2(n6740), .ZN(n7044)
         );
  NAND4_X1 U6129 ( .A1(n7045), .A2(n7046), .A3(n7047), .A4(n7048), .ZN(n3689)
         );
  AOI221_X1 U6130 ( .B1(n6726), .B2(n5275), .C1(n6727), .C2(n5000), .A(n7049), 
        .ZN(n7048) );
  OAI222_X1 U6131 ( .A1(n1082), .A2(n5821), .B1(n1018), .B2(n5828), .C1(n1146), 
        .C2(n5817), .ZN(n7049) );
  AOI221_X1 U6132 ( .B1(n6729), .B2(n5340), .C1(n6730), .C2(n5129), .A(n7050), 
        .ZN(n7047) );
  OAI222_X1 U6133 ( .A1(n570), .A2(n6732), .B1(n506), .B2(n5829), .C1(n762), 
        .C2(n6733), .ZN(n7050) );
  AOI221_X1 U6134 ( .B1(n6734), .B2(n8141), .C1(n6735), .C2(n8077), .A(n7051), 
        .ZN(n7046) );
  OAI222_X1 U6135 ( .A1(n5065), .A2(n6737), .B1(n954), .B2(n5822), .C1(n5468), 
        .C2(n5818), .ZN(n7051) );
  AOI221_X1 U6136 ( .B1(n5832), .B2(DATAIN[39]), .C1(n6738), .C2(OUT1[39]), 
        .A(n7052), .ZN(n7045) );
  OAI22_X1 U6137 ( .A1(n4870), .A2(n5826), .B1(n5404), .B2(n6740), .ZN(n7052)
         );
  NAND4_X1 U6138 ( .A1(n7053), .A2(n7054), .A3(n7055), .A4(n7056), .ZN(n3688)
         );
  AOI221_X1 U6139 ( .B1(n6726), .B2(n5276), .C1(n6727), .C2(n5001), .A(n7057), 
        .ZN(n7056) );
  OAI222_X1 U6140 ( .A1(n1081), .A2(n5821), .B1(n1017), .B2(n5828), .C1(n1145), 
        .C2(n5817), .ZN(n7057) );
  AOI221_X1 U6141 ( .B1(n6729), .B2(n5341), .C1(n6730), .C2(n5130), .A(n7058), 
        .ZN(n7055) );
  OAI222_X1 U6142 ( .A1(n569), .A2(n6732), .B1(n505), .B2(n5829), .C1(n761), 
        .C2(n6733), .ZN(n7058) );
  AOI221_X1 U6143 ( .B1(n6734), .B2(n8140), .C1(n6735), .C2(n8076), .A(n7059), 
        .ZN(n7054) );
  OAI222_X1 U6144 ( .A1(n5066), .A2(n6737), .B1(n953), .B2(n5822), .C1(n5469), 
        .C2(n5818), .ZN(n7059) );
  AOI221_X1 U6145 ( .B1(n5832), .B2(DATAIN[40]), .C1(n6738), .C2(OUT1[40]), 
        .A(n7060), .ZN(n7053) );
  OAI22_X1 U6146 ( .A1(n4871), .A2(n5826), .B1(n5405), .B2(n6740), .ZN(n7060)
         );
  NAND4_X1 U6147 ( .A1(n7061), .A2(n7062), .A3(n7063), .A4(n7064), .ZN(n3687)
         );
  AOI221_X1 U6148 ( .B1(n6726), .B2(n5277), .C1(n6727), .C2(n5002), .A(n7065), 
        .ZN(n7064) );
  OAI222_X1 U6149 ( .A1(n1080), .A2(n5821), .B1(n1016), .B2(n5828), .C1(n1144), 
        .C2(n5817), .ZN(n7065) );
  AOI221_X1 U6150 ( .B1(n6729), .B2(n5342), .C1(n6730), .C2(n5131), .A(n7066), 
        .ZN(n7063) );
  OAI222_X1 U6151 ( .A1(n568), .A2(n6732), .B1(n504), .B2(n5829), .C1(n760), 
        .C2(n6733), .ZN(n7066) );
  AOI221_X1 U6152 ( .B1(n6734), .B2(n8139), .C1(n6735), .C2(n8075), .A(n7067), 
        .ZN(n7062) );
  OAI222_X1 U6153 ( .A1(n5067), .A2(n6737), .B1(n952), .B2(n5822), .C1(n5470), 
        .C2(n5818), .ZN(n7067) );
  AOI221_X1 U6154 ( .B1(n5832), .B2(DATAIN[41]), .C1(n6738), .C2(OUT1[41]), 
        .A(n7068), .ZN(n7061) );
  OAI22_X1 U6155 ( .A1(n4872), .A2(n5826), .B1(n5406), .B2(n6740), .ZN(n7068)
         );
  NAND4_X1 U6156 ( .A1(n7069), .A2(n7070), .A3(n7071), .A4(n7072), .ZN(n3686)
         );
  AOI221_X1 U6157 ( .B1(n6726), .B2(n5278), .C1(n6727), .C2(n5003), .A(n7073), 
        .ZN(n7072) );
  OAI222_X1 U6158 ( .A1(n1079), .A2(n5821), .B1(n1015), .B2(n5828), .C1(n1143), 
        .C2(n5817), .ZN(n7073) );
  AOI221_X1 U6159 ( .B1(n6729), .B2(n5343), .C1(n6730), .C2(n5132), .A(n7074), 
        .ZN(n7071) );
  OAI222_X1 U6160 ( .A1(n567), .A2(n6732), .B1(n503), .B2(n5829), .C1(n759), 
        .C2(n6733), .ZN(n7074) );
  AOI221_X1 U6161 ( .B1(n6734), .B2(n8138), .C1(n6735), .C2(n8074), .A(n7075), 
        .ZN(n7070) );
  OAI222_X1 U6162 ( .A1(n5068), .A2(n6737), .B1(n951), .B2(n5822), .C1(n5471), 
        .C2(n5818), .ZN(n7075) );
  AOI221_X1 U6163 ( .B1(n5832), .B2(DATAIN[42]), .C1(n6738), .C2(OUT1[42]), 
        .A(n7076), .ZN(n7069) );
  OAI22_X1 U6164 ( .A1(n4873), .A2(n5826), .B1(n5407), .B2(n6740), .ZN(n7076)
         );
  NAND4_X1 U6165 ( .A1(n7077), .A2(n7078), .A3(n7079), .A4(n7080), .ZN(n3685)
         );
  AOI221_X1 U6166 ( .B1(n6726), .B2(n5279), .C1(n6727), .C2(n5004), .A(n7081), 
        .ZN(n7080) );
  OAI222_X1 U6167 ( .A1(n1078), .A2(n5821), .B1(n1014), .B2(n5828), .C1(n1142), 
        .C2(n5817), .ZN(n7081) );
  AOI221_X1 U6168 ( .B1(n6729), .B2(n5344), .C1(n6730), .C2(n5133), .A(n7082), 
        .ZN(n7079) );
  OAI222_X1 U6169 ( .A1(n566), .A2(n6732), .B1(n502), .B2(n5829), .C1(n758), 
        .C2(n6733), .ZN(n7082) );
  AOI221_X1 U6170 ( .B1(n6734), .B2(n8137), .C1(n6735), .C2(n8073), .A(n7083), 
        .ZN(n7078) );
  OAI222_X1 U6171 ( .A1(n5069), .A2(n6737), .B1(n950), .B2(n5822), .C1(n5472), 
        .C2(n5818), .ZN(n7083) );
  AOI221_X1 U6172 ( .B1(n5832), .B2(DATAIN[43]), .C1(n6738), .C2(OUT1[43]), 
        .A(n7084), .ZN(n7077) );
  OAI22_X1 U6173 ( .A1(n4874), .A2(n5826), .B1(n5408), .B2(n6740), .ZN(n7084)
         );
  NAND4_X1 U6174 ( .A1(n7085), .A2(n7086), .A3(n7087), .A4(n7088), .ZN(n3684)
         );
  AOI221_X1 U6175 ( .B1(n6726), .B2(n5280), .C1(n6727), .C2(n5005), .A(n7089), 
        .ZN(n7088) );
  OAI222_X1 U6176 ( .A1(n1077), .A2(n5821), .B1(n1013), .B2(n5828), .C1(n1141), 
        .C2(n5817), .ZN(n7089) );
  AOI221_X1 U6177 ( .B1(n6729), .B2(n5345), .C1(n6730), .C2(n5134), .A(n7090), 
        .ZN(n7087) );
  OAI222_X1 U6178 ( .A1(n565), .A2(n6732), .B1(n501), .B2(n5829), .C1(n757), 
        .C2(n6733), .ZN(n7090) );
  AOI221_X1 U6179 ( .B1(n6734), .B2(n8136), .C1(n6735), .C2(n8072), .A(n7091), 
        .ZN(n7086) );
  OAI222_X1 U6180 ( .A1(n5070), .A2(n6737), .B1(n949), .B2(n5822), .C1(n5473), 
        .C2(n5818), .ZN(n7091) );
  AOI221_X1 U6181 ( .B1(n5832), .B2(DATAIN[44]), .C1(n6738), .C2(OUT1[44]), 
        .A(n7092), .ZN(n7085) );
  OAI22_X1 U6182 ( .A1(n4875), .A2(n5826), .B1(n5409), .B2(n6740), .ZN(n7092)
         );
  NAND4_X1 U6183 ( .A1(n7093), .A2(n7094), .A3(n7095), .A4(n7096), .ZN(n3683)
         );
  AOI221_X1 U6184 ( .B1(n6726), .B2(n5281), .C1(n6727), .C2(n5006), .A(n7097), 
        .ZN(n7096) );
  OAI222_X1 U6185 ( .A1(n1076), .A2(n5821), .B1(n1012), .B2(n5828), .C1(n1140), 
        .C2(n5817), .ZN(n7097) );
  AOI221_X1 U6186 ( .B1(n6729), .B2(n5346), .C1(n6730), .C2(n5135), .A(n7098), 
        .ZN(n7095) );
  OAI222_X1 U6187 ( .A1(n564), .A2(n6732), .B1(n500), .B2(n5829), .C1(n756), 
        .C2(n6733), .ZN(n7098) );
  AOI221_X1 U6188 ( .B1(n6734), .B2(n8135), .C1(n6735), .C2(n8071), .A(n7099), 
        .ZN(n7094) );
  OAI222_X1 U6189 ( .A1(n5071), .A2(n6737), .B1(n948), .B2(n5822), .C1(n5474), 
        .C2(n5818), .ZN(n7099) );
  AOI221_X1 U6190 ( .B1(n5832), .B2(DATAIN[45]), .C1(n6738), .C2(OUT1[45]), 
        .A(n7100), .ZN(n7093) );
  OAI22_X1 U6191 ( .A1(n4876), .A2(n5826), .B1(n5410), .B2(n6740), .ZN(n7100)
         );
  NAND4_X1 U6192 ( .A1(n7101), .A2(n7102), .A3(n7103), .A4(n7104), .ZN(n3682)
         );
  AOI221_X1 U6193 ( .B1(n6726), .B2(n5282), .C1(n6727), .C2(n5007), .A(n7105), 
        .ZN(n7104) );
  OAI222_X1 U6194 ( .A1(n1075), .A2(n5821), .B1(n1011), .B2(n5828), .C1(n1139), 
        .C2(n5817), .ZN(n7105) );
  AOI221_X1 U6195 ( .B1(n6729), .B2(n5347), .C1(n6730), .C2(n5136), .A(n7106), 
        .ZN(n7103) );
  OAI222_X1 U6196 ( .A1(n563), .A2(n6732), .B1(n499), .B2(n5829), .C1(n755), 
        .C2(n6733), .ZN(n7106) );
  AOI221_X1 U6197 ( .B1(n6734), .B2(n8134), .C1(n6735), .C2(n8070), .A(n7107), 
        .ZN(n7102) );
  OAI222_X1 U6198 ( .A1(n5072), .A2(n6737), .B1(n947), .B2(n5822), .C1(n5475), 
        .C2(n5818), .ZN(n7107) );
  AOI221_X1 U6199 ( .B1(n5832), .B2(DATAIN[46]), .C1(n6738), .C2(OUT1[46]), 
        .A(n7108), .ZN(n7101) );
  OAI22_X1 U6200 ( .A1(n4877), .A2(n5826), .B1(n5411), .B2(n6740), .ZN(n7108)
         );
  NAND4_X1 U6201 ( .A1(n7109), .A2(n7110), .A3(n7111), .A4(n7112), .ZN(n3681)
         );
  AOI221_X1 U6202 ( .B1(n6726), .B2(n5283), .C1(n6727), .C2(n5008), .A(n7113), 
        .ZN(n7112) );
  OAI222_X1 U6203 ( .A1(n1074), .A2(n5821), .B1(n1010), .B2(n5828), .C1(n1138), 
        .C2(n5817), .ZN(n7113) );
  AOI221_X1 U6204 ( .B1(n6729), .B2(n5348), .C1(n6730), .C2(n5137), .A(n7114), 
        .ZN(n7111) );
  OAI222_X1 U6205 ( .A1(n562), .A2(n6732), .B1(n498), .B2(n5829), .C1(n754), 
        .C2(n6733), .ZN(n7114) );
  AOI221_X1 U6206 ( .B1(n6734), .B2(n8133), .C1(n6735), .C2(n8069), .A(n7115), 
        .ZN(n7110) );
  OAI222_X1 U6207 ( .A1(n5073), .A2(n6737), .B1(n946), .B2(n5822), .C1(n5476), 
        .C2(n5818), .ZN(n7115) );
  AOI221_X1 U6208 ( .B1(n5832), .B2(DATAIN[47]), .C1(n6738), .C2(OUT1[47]), 
        .A(n7116), .ZN(n7109) );
  OAI22_X1 U6209 ( .A1(n4878), .A2(n5826), .B1(n5412), .B2(n6740), .ZN(n7116)
         );
  NAND4_X1 U6210 ( .A1(n7117), .A2(n7118), .A3(n7119), .A4(n7120), .ZN(n3680)
         );
  AOI221_X1 U6211 ( .B1(n6726), .B2(n5284), .C1(n6727), .C2(n5009), .A(n7121), 
        .ZN(n7120) );
  OAI222_X1 U6212 ( .A1(n1073), .A2(n5821), .B1(n1009), .B2(n5828), .C1(n1137), 
        .C2(n5817), .ZN(n7121) );
  AOI221_X1 U6213 ( .B1(n6729), .B2(n5349), .C1(n6730), .C2(n5138), .A(n7122), 
        .ZN(n7119) );
  OAI222_X1 U6214 ( .A1(n561), .A2(n6732), .B1(n497), .B2(n5829), .C1(n753), 
        .C2(n6733), .ZN(n7122) );
  AOI221_X1 U6215 ( .B1(n6734), .B2(n8132), .C1(n6735), .C2(n8068), .A(n7123), 
        .ZN(n7118) );
  OAI222_X1 U6216 ( .A1(n5074), .A2(n6737), .B1(n945), .B2(n5822), .C1(n5477), 
        .C2(n5818), .ZN(n7123) );
  AOI221_X1 U6217 ( .B1(n5832), .B2(DATAIN[48]), .C1(n6738), .C2(OUT1[48]), 
        .A(n7124), .ZN(n7117) );
  OAI22_X1 U6218 ( .A1(n4879), .A2(n5826), .B1(n5413), .B2(n6740), .ZN(n7124)
         );
  NAND4_X1 U6219 ( .A1(n7125), .A2(n7126), .A3(n7127), .A4(n7128), .ZN(n3679)
         );
  AOI221_X1 U6220 ( .B1(n6726), .B2(n5285), .C1(n6727), .C2(n5010), .A(n7129), 
        .ZN(n7128) );
  OAI222_X1 U6221 ( .A1(n1072), .A2(n5821), .B1(n1008), .B2(n5828), .C1(n1136), 
        .C2(n5817), .ZN(n7129) );
  AOI221_X1 U6222 ( .B1(n6729), .B2(n5350), .C1(n6730), .C2(n5139), .A(n7130), 
        .ZN(n7127) );
  OAI222_X1 U6223 ( .A1(n560), .A2(n6732), .B1(n496), .B2(n5829), .C1(n752), 
        .C2(n6733), .ZN(n7130) );
  AOI221_X1 U6224 ( .B1(n6734), .B2(n8131), .C1(n6735), .C2(n8067), .A(n7131), 
        .ZN(n7126) );
  OAI222_X1 U6225 ( .A1(n5075), .A2(n6737), .B1(n944), .B2(n5822), .C1(n5478), 
        .C2(n5818), .ZN(n7131) );
  AOI221_X1 U6226 ( .B1(n5832), .B2(DATAIN[49]), .C1(n6738), .C2(OUT1[49]), 
        .A(n7132), .ZN(n7125) );
  OAI22_X1 U6227 ( .A1(n4880), .A2(n5826), .B1(n5414), .B2(n6740), .ZN(n7132)
         );
  NAND4_X1 U6228 ( .A1(n7133), .A2(n7134), .A3(n7135), .A4(n7136), .ZN(n3678)
         );
  AOI221_X1 U6229 ( .B1(n6726), .B2(n5286), .C1(n6727), .C2(n5011), .A(n7137), 
        .ZN(n7136) );
  OAI222_X1 U6230 ( .A1(n1071), .A2(n5821), .B1(n1007), .B2(n5828), .C1(n1135), 
        .C2(n5817), .ZN(n7137) );
  AOI221_X1 U6231 ( .B1(n6729), .B2(n5351), .C1(n6730), .C2(n5140), .A(n7138), 
        .ZN(n7135) );
  OAI222_X1 U6232 ( .A1(n559), .A2(n6732), .B1(n495), .B2(n5829), .C1(n751), 
        .C2(n6733), .ZN(n7138) );
  AOI221_X1 U6233 ( .B1(n6734), .B2(n8130), .C1(n6735), .C2(n8066), .A(n7139), 
        .ZN(n7134) );
  OAI222_X1 U6234 ( .A1(n5076), .A2(n6737), .B1(n943), .B2(n5822), .C1(n5479), 
        .C2(n5818), .ZN(n7139) );
  AOI221_X1 U6235 ( .B1(n5832), .B2(DATAIN[50]), .C1(n6738), .C2(OUT1[50]), 
        .A(n7140), .ZN(n7133) );
  OAI22_X1 U6236 ( .A1(n4881), .A2(n5826), .B1(n5415), .B2(n6740), .ZN(n7140)
         );
  NAND4_X1 U6237 ( .A1(n7141), .A2(n7142), .A3(n7143), .A4(n7144), .ZN(n3677)
         );
  AOI221_X1 U6238 ( .B1(n6726), .B2(n5287), .C1(n6727), .C2(n5012), .A(n7145), 
        .ZN(n7144) );
  OAI222_X1 U6239 ( .A1(n1070), .A2(n5821), .B1(n1006), .B2(n5828), .C1(n1134), 
        .C2(n5817), .ZN(n7145) );
  AOI221_X1 U6240 ( .B1(n6729), .B2(n5352), .C1(n6730), .C2(n5141), .A(n7146), 
        .ZN(n7143) );
  OAI222_X1 U6241 ( .A1(n558), .A2(n6732), .B1(n494), .B2(n5829), .C1(n750), 
        .C2(n6733), .ZN(n7146) );
  AOI221_X1 U6242 ( .B1(n6734), .B2(n8129), .C1(n6735), .C2(n8065), .A(n7147), 
        .ZN(n7142) );
  OAI222_X1 U6243 ( .A1(n5077), .A2(n6737), .B1(n942), .B2(n5822), .C1(n5480), 
        .C2(n5818), .ZN(n7147) );
  AOI221_X1 U6244 ( .B1(n5832), .B2(DATAIN[51]), .C1(n6738), .C2(OUT1[51]), 
        .A(n7148), .ZN(n7141) );
  OAI22_X1 U6245 ( .A1(n4882), .A2(n5826), .B1(n5416), .B2(n6740), .ZN(n7148)
         );
  NAND4_X1 U6246 ( .A1(n7149), .A2(n7150), .A3(n7151), .A4(n7152), .ZN(n3676)
         );
  AOI221_X1 U6247 ( .B1(n6726), .B2(n5288), .C1(n6727), .C2(n5013), .A(n7153), 
        .ZN(n7152) );
  OAI222_X1 U6248 ( .A1(n1069), .A2(n5821), .B1(n1005), .B2(n5828), .C1(n1133), 
        .C2(n5817), .ZN(n7153) );
  AOI221_X1 U6249 ( .B1(n6729), .B2(n5353), .C1(n6730), .C2(n5142), .A(n7154), 
        .ZN(n7151) );
  OAI222_X1 U6250 ( .A1(n557), .A2(n6732), .B1(n493), .B2(n5829), .C1(n749), 
        .C2(n6733), .ZN(n7154) );
  AOI221_X1 U6251 ( .B1(n6734), .B2(n8128), .C1(n6735), .C2(n8064), .A(n7155), 
        .ZN(n7150) );
  OAI222_X1 U6252 ( .A1(n5078), .A2(n6737), .B1(n941), .B2(n5822), .C1(n5481), 
        .C2(n5818), .ZN(n7155) );
  AOI221_X1 U6253 ( .B1(n5832), .B2(DATAIN[52]), .C1(n6738), .C2(OUT1[52]), 
        .A(n7156), .ZN(n7149) );
  OAI22_X1 U6254 ( .A1(n4883), .A2(n5826), .B1(n5417), .B2(n6740), .ZN(n7156)
         );
  NAND4_X1 U6255 ( .A1(n7157), .A2(n7158), .A3(n7159), .A4(n7160), .ZN(n3675)
         );
  AOI221_X1 U6256 ( .B1(n6726), .B2(n5289), .C1(n6727), .C2(n5014), .A(n7161), 
        .ZN(n7160) );
  OAI222_X1 U6257 ( .A1(n1068), .A2(n5821), .B1(n1004), .B2(n5828), .C1(n1132), 
        .C2(n5817), .ZN(n7161) );
  AOI221_X1 U6258 ( .B1(n6729), .B2(n5354), .C1(n6730), .C2(n5143), .A(n7162), 
        .ZN(n7159) );
  OAI222_X1 U6259 ( .A1(n556), .A2(n6732), .B1(n492), .B2(n5829), .C1(n748), 
        .C2(n6733), .ZN(n7162) );
  AOI221_X1 U6260 ( .B1(n6734), .B2(n8127), .C1(n6735), .C2(n8063), .A(n7163), 
        .ZN(n7158) );
  OAI222_X1 U6261 ( .A1(n5079), .A2(n6737), .B1(n940), .B2(n5822), .C1(n5482), 
        .C2(n5818), .ZN(n7163) );
  AOI221_X1 U6262 ( .B1(n5832), .B2(DATAIN[53]), .C1(n6738), .C2(OUT1[53]), 
        .A(n7164), .ZN(n7157) );
  OAI22_X1 U6263 ( .A1(n4884), .A2(n5826), .B1(n5418), .B2(n6740), .ZN(n7164)
         );
  NAND4_X1 U6264 ( .A1(n7165), .A2(n7166), .A3(n7167), .A4(n7168), .ZN(n3674)
         );
  AOI221_X1 U6265 ( .B1(n6726), .B2(n5290), .C1(n6727), .C2(n5015), .A(n7169), 
        .ZN(n7168) );
  OAI222_X1 U6266 ( .A1(n1067), .A2(n5821), .B1(n1003), .B2(n5828), .C1(n1131), 
        .C2(n5817), .ZN(n7169) );
  AOI221_X1 U6267 ( .B1(n6729), .B2(n5355), .C1(n6730), .C2(n5144), .A(n7170), 
        .ZN(n7167) );
  OAI222_X1 U6268 ( .A1(n555), .A2(n6732), .B1(n491), .B2(n5829), .C1(n747), 
        .C2(n6733), .ZN(n7170) );
  AOI221_X1 U6269 ( .B1(n6734), .B2(n8126), .C1(n6735), .C2(n8062), .A(n7171), 
        .ZN(n7166) );
  OAI222_X1 U6270 ( .A1(n5080), .A2(n6737), .B1(n939), .B2(n5822), .C1(n5483), 
        .C2(n5818), .ZN(n7171) );
  AOI221_X1 U6271 ( .B1(n5832), .B2(DATAIN[54]), .C1(n6738), .C2(OUT1[54]), 
        .A(n7172), .ZN(n7165) );
  OAI22_X1 U6272 ( .A1(n4885), .A2(n5826), .B1(n5419), .B2(n6740), .ZN(n7172)
         );
  NAND4_X1 U6273 ( .A1(n7173), .A2(n7174), .A3(n7175), .A4(n7176), .ZN(n3673)
         );
  AOI221_X1 U6274 ( .B1(n6726), .B2(n5291), .C1(n6727), .C2(n5016), .A(n7177), 
        .ZN(n7176) );
  OAI222_X1 U6275 ( .A1(n1066), .A2(n5821), .B1(n1002), .B2(n5828), .C1(n1130), 
        .C2(n5817), .ZN(n7177) );
  AOI221_X1 U6276 ( .B1(n6729), .B2(n5356), .C1(n6730), .C2(n5145), .A(n7178), 
        .ZN(n7175) );
  OAI222_X1 U6277 ( .A1(n554), .A2(n6732), .B1(n490), .B2(n5829), .C1(n746), 
        .C2(n6733), .ZN(n7178) );
  AOI221_X1 U6278 ( .B1(n6734), .B2(n8125), .C1(n6735), .C2(n8061), .A(n7179), 
        .ZN(n7174) );
  OAI222_X1 U6279 ( .A1(n5081), .A2(n6737), .B1(n938), .B2(n5822), .C1(n5484), 
        .C2(n5818), .ZN(n7179) );
  AOI221_X1 U6280 ( .B1(n5832), .B2(DATAIN[55]), .C1(n6738), .C2(OUT1[55]), 
        .A(n7180), .ZN(n7173) );
  OAI22_X1 U6281 ( .A1(n4886), .A2(n5826), .B1(n5420), .B2(n6740), .ZN(n7180)
         );
  NAND4_X1 U6282 ( .A1(n7181), .A2(n7182), .A3(n7183), .A4(n7184), .ZN(n3672)
         );
  AOI221_X1 U6283 ( .B1(n6726), .B2(n5292), .C1(n6727), .C2(n5017), .A(n7185), 
        .ZN(n7184) );
  OAI222_X1 U6284 ( .A1(n1065), .A2(n5821), .B1(n1001), .B2(n5828), .C1(n1129), 
        .C2(n5817), .ZN(n7185) );
  AOI221_X1 U6285 ( .B1(n6729), .B2(n5357), .C1(n6730), .C2(n5146), .A(n7186), 
        .ZN(n7183) );
  OAI222_X1 U6286 ( .A1(n553), .A2(n6732), .B1(n489), .B2(n5829), .C1(n745), 
        .C2(n6733), .ZN(n7186) );
  AOI221_X1 U6287 ( .B1(n6734), .B2(n8124), .C1(n6735), .C2(n8060), .A(n7187), 
        .ZN(n7182) );
  OAI222_X1 U6288 ( .A1(n5082), .A2(n6737), .B1(n937), .B2(n5822), .C1(n5485), 
        .C2(n5818), .ZN(n7187) );
  AOI221_X1 U6289 ( .B1(n5832), .B2(DATAIN[56]), .C1(n6738), .C2(OUT1[56]), 
        .A(n7188), .ZN(n7181) );
  OAI22_X1 U6290 ( .A1(n4887), .A2(n5826), .B1(n5421), .B2(n6740), .ZN(n7188)
         );
  NAND4_X1 U6291 ( .A1(n7189), .A2(n7190), .A3(n7191), .A4(n7192), .ZN(n3671)
         );
  AOI221_X1 U6292 ( .B1(n6726), .B2(n5293), .C1(n6727), .C2(n5018), .A(n7193), 
        .ZN(n7192) );
  OAI222_X1 U6293 ( .A1(n1064), .A2(n5821), .B1(n1000), .B2(n5828), .C1(n1128), 
        .C2(n5817), .ZN(n7193) );
  AOI221_X1 U6294 ( .B1(n6729), .B2(n5358), .C1(n6730), .C2(n5147), .A(n7194), 
        .ZN(n7191) );
  OAI222_X1 U6295 ( .A1(n552), .A2(n6732), .B1(n488), .B2(n5829), .C1(n744), 
        .C2(n6733), .ZN(n7194) );
  AOI221_X1 U6296 ( .B1(n6734), .B2(n8123), .C1(n6735), .C2(n8059), .A(n7195), 
        .ZN(n7190) );
  OAI222_X1 U6297 ( .A1(n5083), .A2(n6737), .B1(n936), .B2(n5822), .C1(n5486), 
        .C2(n5818), .ZN(n7195) );
  AOI221_X1 U6298 ( .B1(n5832), .B2(DATAIN[57]), .C1(n6738), .C2(OUT1[57]), 
        .A(n7196), .ZN(n7189) );
  OAI22_X1 U6299 ( .A1(n4888), .A2(n5826), .B1(n5422), .B2(n6740), .ZN(n7196)
         );
  NAND4_X1 U6300 ( .A1(n7197), .A2(n7198), .A3(n7199), .A4(n7200), .ZN(n3670)
         );
  AOI221_X1 U6301 ( .B1(n6726), .B2(n5294), .C1(n6727), .C2(n5019), .A(n7201), 
        .ZN(n7200) );
  OAI222_X1 U6302 ( .A1(n1063), .A2(n5821), .B1(n999), .B2(n5828), .C1(n1127), 
        .C2(n5817), .ZN(n7201) );
  AOI221_X1 U6303 ( .B1(n6729), .B2(n5359), .C1(n6730), .C2(n5148), .A(n7202), 
        .ZN(n7199) );
  OAI222_X1 U6304 ( .A1(n551), .A2(n6732), .B1(n487), .B2(n5829), .C1(n743), 
        .C2(n6733), .ZN(n7202) );
  AOI221_X1 U6305 ( .B1(n6734), .B2(n8122), .C1(n6735), .C2(n8058), .A(n7203), 
        .ZN(n7198) );
  OAI222_X1 U6306 ( .A1(n5084), .A2(n6737), .B1(n935), .B2(n5822), .C1(n5487), 
        .C2(n5818), .ZN(n7203) );
  AOI221_X1 U6307 ( .B1(n5832), .B2(DATAIN[58]), .C1(n6738), .C2(OUT1[58]), 
        .A(n7204), .ZN(n7197) );
  OAI22_X1 U6308 ( .A1(n4889), .A2(n5826), .B1(n5423), .B2(n6740), .ZN(n7204)
         );
  NAND4_X1 U6309 ( .A1(n7205), .A2(n7206), .A3(n7207), .A4(n7208), .ZN(n3669)
         );
  AOI221_X1 U6310 ( .B1(n6726), .B2(n5295), .C1(n6727), .C2(n5020), .A(n7209), 
        .ZN(n7208) );
  OAI222_X1 U6311 ( .A1(n1062), .A2(n5821), .B1(n998), .B2(n5828), .C1(n1126), 
        .C2(n5817), .ZN(n7209) );
  AOI221_X1 U6312 ( .B1(n6729), .B2(n5360), .C1(n6730), .C2(n5149), .A(n7210), 
        .ZN(n7207) );
  OAI222_X1 U6313 ( .A1(n550), .A2(n6732), .B1(n486), .B2(n5829), .C1(n742), 
        .C2(n6733), .ZN(n7210) );
  AOI221_X1 U6314 ( .B1(n6734), .B2(n8121), .C1(n6735), .C2(n8057), .A(n7211), 
        .ZN(n7206) );
  OAI222_X1 U6315 ( .A1(n5085), .A2(n6737), .B1(n934), .B2(n5822), .C1(n5488), 
        .C2(n5818), .ZN(n7211) );
  AOI221_X1 U6316 ( .B1(n5832), .B2(DATAIN[59]), .C1(n6738), .C2(OUT1[59]), 
        .A(n7212), .ZN(n7205) );
  OAI22_X1 U6317 ( .A1(n4890), .A2(n5826), .B1(n5424), .B2(n6740), .ZN(n7212)
         );
  NAND4_X1 U6318 ( .A1(n7213), .A2(n7214), .A3(n7215), .A4(n7216), .ZN(n3668)
         );
  AOI221_X1 U6319 ( .B1(n6726), .B2(n5296), .C1(n6727), .C2(n5021), .A(n7217), 
        .ZN(n7216) );
  OAI222_X1 U6320 ( .A1(n1061), .A2(n5821), .B1(n997), .B2(n5828), .C1(n1125), 
        .C2(n5817), .ZN(n7217) );
  AOI221_X1 U6321 ( .B1(n6729), .B2(n5361), .C1(n6730), .C2(n5150), .A(n7218), 
        .ZN(n7215) );
  OAI222_X1 U6322 ( .A1(n549), .A2(n6732), .B1(n485), .B2(n5829), .C1(n741), 
        .C2(n6733), .ZN(n7218) );
  AOI221_X1 U6323 ( .B1(n6734), .B2(n8120), .C1(n6735), .C2(n8056), .A(n7219), 
        .ZN(n7214) );
  OAI222_X1 U6324 ( .A1(n5086), .A2(n6737), .B1(n933), .B2(n5822), .C1(n5489), 
        .C2(n5818), .ZN(n7219) );
  AOI221_X1 U6325 ( .B1(n5832), .B2(DATAIN[60]), .C1(n6738), .C2(OUT1[60]), 
        .A(n7220), .ZN(n7213) );
  OAI22_X1 U6326 ( .A1(n4891), .A2(n5826), .B1(n5425), .B2(n6740), .ZN(n7220)
         );
  NAND4_X1 U6327 ( .A1(n7221), .A2(n7222), .A3(n7223), .A4(n7224), .ZN(n3667)
         );
  AOI221_X1 U6328 ( .B1(n6726), .B2(n5297), .C1(n6727), .C2(n5022), .A(n7225), 
        .ZN(n7224) );
  OAI222_X1 U6329 ( .A1(n1060), .A2(n5821), .B1(n996), .B2(n5828), .C1(n1124), 
        .C2(n5817), .ZN(n7225) );
  AOI221_X1 U6330 ( .B1(n6729), .B2(n5362), .C1(n6730), .C2(n5151), .A(n7226), 
        .ZN(n7223) );
  OAI222_X1 U6331 ( .A1(n548), .A2(n6732), .B1(n484), .B2(n5829), .C1(n740), 
        .C2(n6733), .ZN(n7226) );
  AOI221_X1 U6332 ( .B1(n6734), .B2(n8119), .C1(n6735), .C2(n8055), .A(n7227), 
        .ZN(n7222) );
  OAI222_X1 U6333 ( .A1(n5087), .A2(n6737), .B1(n932), .B2(n5822), .C1(n5490), 
        .C2(n5818), .ZN(n7227) );
  AOI221_X1 U6334 ( .B1(n5832), .B2(DATAIN[61]), .C1(n6738), .C2(OUT1[61]), 
        .A(n7228), .ZN(n7221) );
  OAI22_X1 U6335 ( .A1(n4892), .A2(n5826), .B1(n5426), .B2(n6740), .ZN(n7228)
         );
  NAND4_X1 U6336 ( .A1(n7229), .A2(n7230), .A3(n7231), .A4(n7232), .ZN(n3666)
         );
  AOI221_X1 U6337 ( .B1(n6726), .B2(n5298), .C1(n6727), .C2(n5023), .A(n7233), 
        .ZN(n7232) );
  OAI222_X1 U6338 ( .A1(n1059), .A2(n5821), .B1(n995), .B2(n5828), .C1(n1123), 
        .C2(n5817), .ZN(n7233) );
  AOI221_X1 U6339 ( .B1(n6729), .B2(n5363), .C1(n6730), .C2(n5152), .A(n7234), 
        .ZN(n7231) );
  OAI222_X1 U6340 ( .A1(n547), .A2(n6732), .B1(n483), .B2(n5829), .C1(n739), 
        .C2(n6733), .ZN(n7234) );
  AOI221_X1 U6341 ( .B1(n6734), .B2(n8118), .C1(n6735), .C2(n8054), .A(n7235), 
        .ZN(n7230) );
  OAI222_X1 U6342 ( .A1(n5088), .A2(n6737), .B1(n931), .B2(n5822), .C1(n5491), 
        .C2(n5818), .ZN(n7235) );
  AOI221_X1 U6343 ( .B1(n5832), .B2(DATAIN[62]), .C1(n6738), .C2(OUT1[62]), 
        .A(n7236), .ZN(n7229) );
  OAI22_X1 U6344 ( .A1(n4893), .A2(n5826), .B1(n5427), .B2(n6740), .ZN(n7236)
         );
  NAND4_X1 U6345 ( .A1(n7237), .A2(n7238), .A3(n7239), .A4(n7240), .ZN(n3665)
         );
  AOI221_X1 U6346 ( .B1(n6726), .B2(n5299), .C1(n6727), .C2(n5024), .A(n7241), 
        .ZN(n7240) );
  OAI222_X1 U6347 ( .A1(n1058), .A2(n5821), .B1(n994), .B2(n5828), .C1(n1122), 
        .C2(n5817), .ZN(n7241) );
  AND3_X1 U6348 ( .A1(N333), .A2(n5851), .A3(N334), .ZN(n7242) );
  AOI221_X1 U6349 ( .B1(n6729), .B2(n5364), .C1(n6730), .C2(n5153), .A(n7250), 
        .ZN(n7239) );
  OAI222_X1 U6350 ( .A1(n546), .A2(n6732), .B1(n482), .B2(n5829), .C1(n738), 
        .C2(n6733), .ZN(n7250) );
  NOR3_X1 U6351 ( .A1(N332), .A2(N333), .A3(n5867), .ZN(n7249) );
  NOR2_X1 U6352 ( .A1(n7244), .A2(n5851), .ZN(n7246) );
  AOI221_X1 U6353 ( .B1(n6734), .B2(n8117), .C1(n6735), .C2(n8053), .A(n7253), 
        .ZN(n7238) );
  OAI222_X1 U6354 ( .A1(n5089), .A2(n6737), .B1(n930), .B2(n5822), .C1(n5492), 
        .C2(n5818), .ZN(n7253) );
  AND2_X1 U6355 ( .A1(n7243), .A2(N334), .ZN(n7245) );
  INV_X1 U6356 ( .A(n7255), .ZN(n7243) );
  AND2_X1 U6357 ( .A1(n7248), .A2(N333), .ZN(n7251) );
  AOI221_X1 U6358 ( .B1(n5832), .B2(DATAIN[63]), .C1(n6738), .C2(OUT1[63]), 
        .A(n7256), .ZN(n7237) );
  OAI22_X1 U6359 ( .A1(n4894), .A2(n5826), .B1(n5428), .B2(n6740), .ZN(n7256)
         );
  NOR3_X1 U6360 ( .A1(n5867), .A2(N333), .A3(n7244), .ZN(n7252) );
  INV_X1 U6361 ( .A(N332), .ZN(n7244) );
  INV_X1 U6362 ( .A(n5856), .ZN(n7257) );
  INV_X1 U6363 ( .A(N333), .ZN(n7247) );
  NOR2_X1 U6364 ( .A1(n7255), .A2(N334), .ZN(n7248) );
  NAND3_X1 U6365 ( .A1(n7258), .A2(n6455), .A3(n7259), .ZN(n7255) );
  NOR2_X1 U6366 ( .A1(N332), .A2(n5851), .ZN(n7254) );
  NAND4_X1 U6367 ( .A1(n7260), .A2(n7261), .A3(WR), .A4(n7262), .ZN(n7259) );
  NOR3_X1 U6368 ( .A1(n7263), .A2(n7264), .A3(n7265), .ZN(n7262) );
  XOR2_X1 U6369 ( .A(n6631), .B(N557), .Z(n7264) );
  XNOR2_X1 U6370 ( .A(N556), .B(n6644), .ZN(n7261) );
  XOR2_X1 U6371 ( .A(N555), .B(n6643), .Z(n7260) );
  NAND2_X1 U6372 ( .A1(n7266), .A2(n6455), .ZN(n7258) );
  NAND4_X1 U6373 ( .A1(n7267), .A2(n7268), .A3(n7269), .A4(n7270), .ZN(n3664)
         );
  AOI221_X1 U6374 ( .B1(n7271), .B2(n5236), .C1(n7272), .C2(n4961), .A(n7273), 
        .ZN(n7270) );
  OAI222_X1 U6375 ( .A1(n1121), .A2(n5820), .B1(n1057), .B2(n5823), .C1(n1185), 
        .C2(n5815), .ZN(n7273) );
  AOI221_X1 U6376 ( .B1(n7274), .B2(n5301), .C1(n7275), .C2(n5090), .A(n7276), 
        .ZN(n7269) );
  OAI222_X1 U6377 ( .A1(n609), .A2(n7277), .B1(n545), .B2(n5824), .C1(n801), 
        .C2(n7278), .ZN(n7276) );
  AOI221_X1 U6378 ( .B1(n7279), .B2(n8180), .C1(n7280), .C2(n8116), .A(n7281), 
        .ZN(n7268) );
  OAI222_X1 U6379 ( .A1(n5026), .A2(n7282), .B1(n993), .B2(n5825), .C1(n5429), 
        .C2(n5816), .ZN(n7281) );
  AOI221_X1 U6380 ( .B1(n5833), .B2(DATAIN[0]), .C1(n7283), .C2(OUT2[0]), .A(
        n7284), .ZN(n7267) );
  OAI22_X1 U6381 ( .A1(n4831), .A2(n5827), .B1(n5365), .B2(n7285), .ZN(n7284)
         );
  NAND4_X1 U6382 ( .A1(n7286), .A2(n7287), .A3(n7288), .A4(n7289), .ZN(n3663)
         );
  AOI221_X1 U6383 ( .B1(n7271), .B2(n5237), .C1(n7272), .C2(n4962), .A(n7290), 
        .ZN(n7289) );
  OAI222_X1 U6384 ( .A1(n1120), .A2(n5820), .B1(n1056), .B2(n5823), .C1(n1184), 
        .C2(n5815), .ZN(n7290) );
  AOI221_X1 U6385 ( .B1(n7274), .B2(n5302), .C1(n7275), .C2(n5091), .A(n7291), 
        .ZN(n7288) );
  OAI222_X1 U6386 ( .A1(n608), .A2(n7277), .B1(n544), .B2(n5824), .C1(n800), 
        .C2(n7278), .ZN(n7291) );
  AOI221_X1 U6387 ( .B1(n7279), .B2(n8179), .C1(n7280), .C2(n8115), .A(n7292), 
        .ZN(n7287) );
  OAI222_X1 U6388 ( .A1(n5027), .A2(n7282), .B1(n992), .B2(n5825), .C1(n5430), 
        .C2(n5816), .ZN(n7292) );
  AOI221_X1 U6389 ( .B1(n5833), .B2(DATAIN[1]), .C1(n7283), .C2(OUT2[1]), .A(
        n7293), .ZN(n7286) );
  OAI22_X1 U6390 ( .A1(n4832), .A2(n5827), .B1(n5366), .B2(n7285), .ZN(n7293)
         );
  NAND4_X1 U6391 ( .A1(n7294), .A2(n7295), .A3(n7296), .A4(n7297), .ZN(n3662)
         );
  AOI221_X1 U6392 ( .B1(n7271), .B2(n5238), .C1(n7272), .C2(n4963), .A(n7298), 
        .ZN(n7297) );
  OAI222_X1 U6393 ( .A1(n1119), .A2(n5820), .B1(n1055), .B2(n5823), .C1(n1183), 
        .C2(n5815), .ZN(n7298) );
  AOI221_X1 U6394 ( .B1(n7274), .B2(n5303), .C1(n7275), .C2(n5092), .A(n7299), 
        .ZN(n7296) );
  OAI222_X1 U6395 ( .A1(n607), .A2(n7277), .B1(n543), .B2(n5824), .C1(n799), 
        .C2(n7278), .ZN(n7299) );
  AOI221_X1 U6396 ( .B1(n7279), .B2(n8178), .C1(n7280), .C2(n8114), .A(n7300), 
        .ZN(n7295) );
  OAI222_X1 U6397 ( .A1(n5028), .A2(n7282), .B1(n991), .B2(n5825), .C1(n5431), 
        .C2(n5816), .ZN(n7300) );
  AOI221_X1 U6398 ( .B1(n5833), .B2(DATAIN[2]), .C1(n7283), .C2(OUT2[2]), .A(
        n7301), .ZN(n7294) );
  OAI22_X1 U6399 ( .A1(n4833), .A2(n5827), .B1(n5367), .B2(n7285), .ZN(n7301)
         );
  NAND4_X1 U6400 ( .A1(n7302), .A2(n7303), .A3(n7304), .A4(n7305), .ZN(n3661)
         );
  AOI221_X1 U6401 ( .B1(n7271), .B2(n5239), .C1(n7272), .C2(n4964), .A(n7306), 
        .ZN(n7305) );
  OAI222_X1 U6402 ( .A1(n1118), .A2(n5820), .B1(n1054), .B2(n5823), .C1(n1182), 
        .C2(n5815), .ZN(n7306) );
  AOI221_X1 U6403 ( .B1(n7274), .B2(n5304), .C1(n7275), .C2(n5093), .A(n7307), 
        .ZN(n7304) );
  OAI222_X1 U6404 ( .A1(n606), .A2(n7277), .B1(n542), .B2(n5824), .C1(n798), 
        .C2(n7278), .ZN(n7307) );
  AOI221_X1 U6405 ( .B1(n7279), .B2(n8177), .C1(n7280), .C2(n8113), .A(n7308), 
        .ZN(n7303) );
  OAI222_X1 U6406 ( .A1(n5029), .A2(n7282), .B1(n990), .B2(n5825), .C1(n5432), 
        .C2(n5816), .ZN(n7308) );
  AOI221_X1 U6407 ( .B1(n5833), .B2(DATAIN[3]), .C1(n7283), .C2(OUT2[3]), .A(
        n7309), .ZN(n7302) );
  OAI22_X1 U6408 ( .A1(n4834), .A2(n5827), .B1(n5368), .B2(n7285), .ZN(n7309)
         );
  NAND4_X1 U6409 ( .A1(n7310), .A2(n7311), .A3(n7312), .A4(n7313), .ZN(n3660)
         );
  AOI221_X1 U6410 ( .B1(n7271), .B2(n5240), .C1(n7272), .C2(n4965), .A(n7314), 
        .ZN(n7313) );
  OAI222_X1 U6411 ( .A1(n1117), .A2(n5820), .B1(n1053), .B2(n5823), .C1(n1181), 
        .C2(n5815), .ZN(n7314) );
  AOI221_X1 U6412 ( .B1(n7274), .B2(n5305), .C1(n7275), .C2(n5094), .A(n7315), 
        .ZN(n7312) );
  OAI222_X1 U6413 ( .A1(n605), .A2(n7277), .B1(n541), .B2(n5824), .C1(n797), 
        .C2(n7278), .ZN(n7315) );
  AOI221_X1 U6414 ( .B1(n7279), .B2(n8176), .C1(n7280), .C2(n8112), .A(n7316), 
        .ZN(n7311) );
  OAI222_X1 U6415 ( .A1(n5030), .A2(n7282), .B1(n989), .B2(n5825), .C1(n5433), 
        .C2(n5816), .ZN(n7316) );
  AOI221_X1 U6416 ( .B1(n5833), .B2(DATAIN[4]), .C1(n7283), .C2(OUT2[4]), .A(
        n7317), .ZN(n7310) );
  OAI22_X1 U6417 ( .A1(n4835), .A2(n5827), .B1(n5369), .B2(n7285), .ZN(n7317)
         );
  NAND4_X1 U6418 ( .A1(n7318), .A2(n7319), .A3(n7320), .A4(n7321), .ZN(n3659)
         );
  AOI221_X1 U6419 ( .B1(n7271), .B2(n5241), .C1(n7272), .C2(n4966), .A(n7322), 
        .ZN(n7321) );
  OAI222_X1 U6420 ( .A1(n1116), .A2(n5820), .B1(n1052), .B2(n5823), .C1(n1180), 
        .C2(n5815), .ZN(n7322) );
  AOI221_X1 U6421 ( .B1(n7274), .B2(n5306), .C1(n7275), .C2(n5095), .A(n7323), 
        .ZN(n7320) );
  OAI222_X1 U6422 ( .A1(n604), .A2(n7277), .B1(n540), .B2(n5824), .C1(n796), 
        .C2(n7278), .ZN(n7323) );
  AOI221_X1 U6423 ( .B1(n7279), .B2(n8175), .C1(n7280), .C2(n8111), .A(n7324), 
        .ZN(n7319) );
  OAI222_X1 U6424 ( .A1(n5031), .A2(n7282), .B1(n988), .B2(n5825), .C1(n5434), 
        .C2(n5816), .ZN(n7324) );
  AOI221_X1 U6425 ( .B1(n5833), .B2(DATAIN[5]), .C1(n7283), .C2(OUT2[5]), .A(
        n7325), .ZN(n7318) );
  OAI22_X1 U6426 ( .A1(n4836), .A2(n5827), .B1(n5370), .B2(n7285), .ZN(n7325)
         );
  NAND4_X1 U6427 ( .A1(n7326), .A2(n7327), .A3(n7328), .A4(n7329), .ZN(n3658)
         );
  AOI221_X1 U6428 ( .B1(n7271), .B2(n5242), .C1(n7272), .C2(n4967), .A(n7330), 
        .ZN(n7329) );
  OAI222_X1 U6429 ( .A1(n1115), .A2(n5820), .B1(n1051), .B2(n5823), .C1(n1179), 
        .C2(n5815), .ZN(n7330) );
  AOI221_X1 U6430 ( .B1(n7274), .B2(n5307), .C1(n7275), .C2(n5096), .A(n7331), 
        .ZN(n7328) );
  OAI222_X1 U6431 ( .A1(n603), .A2(n7277), .B1(n539), .B2(n5824), .C1(n795), 
        .C2(n7278), .ZN(n7331) );
  AOI221_X1 U6432 ( .B1(n7279), .B2(n8174), .C1(n7280), .C2(n8110), .A(n7332), 
        .ZN(n7327) );
  OAI222_X1 U6433 ( .A1(n5032), .A2(n7282), .B1(n987), .B2(n5825), .C1(n5435), 
        .C2(n5816), .ZN(n7332) );
  AOI221_X1 U6434 ( .B1(n5833), .B2(DATAIN[6]), .C1(n7283), .C2(OUT2[6]), .A(
        n7333), .ZN(n7326) );
  OAI22_X1 U6435 ( .A1(n4837), .A2(n5827), .B1(n5371), .B2(n7285), .ZN(n7333)
         );
  NAND4_X1 U6436 ( .A1(n7334), .A2(n7335), .A3(n7336), .A4(n7337), .ZN(n3657)
         );
  AOI221_X1 U6437 ( .B1(n7271), .B2(n5243), .C1(n7272), .C2(n4968), .A(n7338), 
        .ZN(n7337) );
  OAI222_X1 U6438 ( .A1(n1114), .A2(n5820), .B1(n1050), .B2(n5823), .C1(n1178), 
        .C2(n5815), .ZN(n7338) );
  AOI221_X1 U6439 ( .B1(n7274), .B2(n5308), .C1(n7275), .C2(n5097), .A(n7339), 
        .ZN(n7336) );
  OAI222_X1 U6440 ( .A1(n602), .A2(n7277), .B1(n538), .B2(n5824), .C1(n794), 
        .C2(n7278), .ZN(n7339) );
  AOI221_X1 U6441 ( .B1(n7279), .B2(n8173), .C1(n7280), .C2(n8109), .A(n7340), 
        .ZN(n7335) );
  OAI222_X1 U6442 ( .A1(n5033), .A2(n7282), .B1(n986), .B2(n5825), .C1(n5436), 
        .C2(n5816), .ZN(n7340) );
  AOI221_X1 U6443 ( .B1(n5833), .B2(DATAIN[7]), .C1(n7283), .C2(OUT2[7]), .A(
        n7341), .ZN(n7334) );
  OAI22_X1 U6444 ( .A1(n4838), .A2(n5827), .B1(n5372), .B2(n7285), .ZN(n7341)
         );
  NAND4_X1 U6445 ( .A1(n7342), .A2(n7343), .A3(n7344), .A4(n7345), .ZN(n3656)
         );
  AOI221_X1 U6446 ( .B1(n7271), .B2(n5244), .C1(n7272), .C2(n4969), .A(n7346), 
        .ZN(n7345) );
  OAI222_X1 U6447 ( .A1(n1113), .A2(n5820), .B1(n1049), .B2(n5823), .C1(n1177), 
        .C2(n5815), .ZN(n7346) );
  AOI221_X1 U6448 ( .B1(n7274), .B2(n5309), .C1(n7275), .C2(n5098), .A(n7347), 
        .ZN(n7344) );
  OAI222_X1 U6449 ( .A1(n601), .A2(n7277), .B1(n537), .B2(n5824), .C1(n793), 
        .C2(n7278), .ZN(n7347) );
  AOI221_X1 U6450 ( .B1(n7279), .B2(n8172), .C1(n7280), .C2(n8108), .A(n7348), 
        .ZN(n7343) );
  OAI222_X1 U6451 ( .A1(n5034), .A2(n7282), .B1(n985), .B2(n5825), .C1(n5437), 
        .C2(n5816), .ZN(n7348) );
  AOI221_X1 U6452 ( .B1(n5833), .B2(DATAIN[8]), .C1(n7283), .C2(OUT2[8]), .A(
        n7349), .ZN(n7342) );
  OAI22_X1 U6453 ( .A1(n4839), .A2(n5827), .B1(n5373), .B2(n7285), .ZN(n7349)
         );
  NAND4_X1 U6454 ( .A1(n7350), .A2(n7351), .A3(n7352), .A4(n7353), .ZN(n3655)
         );
  AOI221_X1 U6455 ( .B1(n7271), .B2(n5245), .C1(n7272), .C2(n4970), .A(n7354), 
        .ZN(n7353) );
  OAI222_X1 U6456 ( .A1(n1112), .A2(n5820), .B1(n1048), .B2(n5823), .C1(n1176), 
        .C2(n5815), .ZN(n7354) );
  AOI221_X1 U6457 ( .B1(n7274), .B2(n5310), .C1(n7275), .C2(n5099), .A(n7355), 
        .ZN(n7352) );
  OAI222_X1 U6458 ( .A1(n600), .A2(n7277), .B1(n536), .B2(n5824), .C1(n792), 
        .C2(n7278), .ZN(n7355) );
  AOI221_X1 U6459 ( .B1(n7279), .B2(n8171), .C1(n7280), .C2(n8107), .A(n7356), 
        .ZN(n7351) );
  OAI222_X1 U6460 ( .A1(n5035), .A2(n7282), .B1(n984), .B2(n5825), .C1(n5438), 
        .C2(n5816), .ZN(n7356) );
  AOI221_X1 U6461 ( .B1(n5833), .B2(DATAIN[9]), .C1(n7283), .C2(OUT2[9]), .A(
        n7357), .ZN(n7350) );
  OAI22_X1 U6462 ( .A1(n4840), .A2(n5827), .B1(n5374), .B2(n7285), .ZN(n7357)
         );
  NAND4_X1 U6463 ( .A1(n7358), .A2(n7359), .A3(n7360), .A4(n7361), .ZN(n3654)
         );
  AOI221_X1 U6464 ( .B1(n7271), .B2(n5246), .C1(n7272), .C2(n4971), .A(n7362), 
        .ZN(n7361) );
  OAI222_X1 U6465 ( .A1(n1111), .A2(n5820), .B1(n1047), .B2(n5823), .C1(n1175), 
        .C2(n5815), .ZN(n7362) );
  AOI221_X1 U6466 ( .B1(n7274), .B2(n5311), .C1(n7275), .C2(n5100), .A(n7363), 
        .ZN(n7360) );
  OAI222_X1 U6467 ( .A1(n599), .A2(n7277), .B1(n535), .B2(n5824), .C1(n791), 
        .C2(n7278), .ZN(n7363) );
  AOI221_X1 U6468 ( .B1(n7279), .B2(n8170), .C1(n7280), .C2(n8106), .A(n7364), 
        .ZN(n7359) );
  OAI222_X1 U6469 ( .A1(n5036), .A2(n7282), .B1(n983), .B2(n5825), .C1(n5439), 
        .C2(n5816), .ZN(n7364) );
  AOI221_X1 U6470 ( .B1(n5833), .B2(DATAIN[10]), .C1(n7283), .C2(OUT2[10]), 
        .A(n7365), .ZN(n7358) );
  OAI22_X1 U6471 ( .A1(n4841), .A2(n5827), .B1(n5375), .B2(n7285), .ZN(n7365)
         );
  NAND4_X1 U6472 ( .A1(n7366), .A2(n7367), .A3(n7368), .A4(n7369), .ZN(n3653)
         );
  AOI221_X1 U6473 ( .B1(n7271), .B2(n5247), .C1(n7272), .C2(n4972), .A(n7370), 
        .ZN(n7369) );
  OAI222_X1 U6474 ( .A1(n1110), .A2(n5820), .B1(n1046), .B2(n5823), .C1(n1174), 
        .C2(n5815), .ZN(n7370) );
  AOI221_X1 U6475 ( .B1(n7274), .B2(n5312), .C1(n7275), .C2(n5101), .A(n7371), 
        .ZN(n7368) );
  OAI222_X1 U6476 ( .A1(n598), .A2(n7277), .B1(n534), .B2(n5824), .C1(n790), 
        .C2(n7278), .ZN(n7371) );
  AOI221_X1 U6477 ( .B1(n7279), .B2(n8169), .C1(n7280), .C2(n8105), .A(n7372), 
        .ZN(n7367) );
  OAI222_X1 U6478 ( .A1(n5037), .A2(n7282), .B1(n982), .B2(n5825), .C1(n5440), 
        .C2(n5816), .ZN(n7372) );
  AOI221_X1 U6479 ( .B1(n5833), .B2(DATAIN[11]), .C1(n7283), .C2(OUT2[11]), 
        .A(n7373), .ZN(n7366) );
  OAI22_X1 U6480 ( .A1(n4842), .A2(n5827), .B1(n5376), .B2(n7285), .ZN(n7373)
         );
  NAND4_X1 U6481 ( .A1(n7374), .A2(n7375), .A3(n7376), .A4(n7377), .ZN(n3652)
         );
  AOI221_X1 U6482 ( .B1(n7271), .B2(n5248), .C1(n7272), .C2(n4973), .A(n7378), 
        .ZN(n7377) );
  OAI222_X1 U6483 ( .A1(n1109), .A2(n5820), .B1(n1045), .B2(n5823), .C1(n1173), 
        .C2(n5815), .ZN(n7378) );
  AOI221_X1 U6484 ( .B1(n7274), .B2(n5313), .C1(n7275), .C2(n5102), .A(n7379), 
        .ZN(n7376) );
  OAI222_X1 U6485 ( .A1(n597), .A2(n7277), .B1(n533), .B2(n5824), .C1(n789), 
        .C2(n7278), .ZN(n7379) );
  AOI221_X1 U6486 ( .B1(n7279), .B2(n8168), .C1(n7280), .C2(n8104), .A(n7380), 
        .ZN(n7375) );
  OAI222_X1 U6487 ( .A1(n5038), .A2(n7282), .B1(n981), .B2(n5825), .C1(n5441), 
        .C2(n5816), .ZN(n7380) );
  AOI221_X1 U6488 ( .B1(n5833), .B2(DATAIN[12]), .C1(n7283), .C2(OUT2[12]), 
        .A(n7381), .ZN(n7374) );
  OAI22_X1 U6489 ( .A1(n4843), .A2(n5827), .B1(n5377), .B2(n7285), .ZN(n7381)
         );
  NAND4_X1 U6490 ( .A1(n7382), .A2(n7383), .A3(n7384), .A4(n7385), .ZN(n3651)
         );
  AOI221_X1 U6491 ( .B1(n7271), .B2(n5249), .C1(n7272), .C2(n4974), .A(n7386), 
        .ZN(n7385) );
  OAI222_X1 U6492 ( .A1(n1108), .A2(n5820), .B1(n1044), .B2(n5823), .C1(n1172), 
        .C2(n5815), .ZN(n7386) );
  AOI221_X1 U6493 ( .B1(n7274), .B2(n5314), .C1(n7275), .C2(n5103), .A(n7387), 
        .ZN(n7384) );
  OAI222_X1 U6494 ( .A1(n596), .A2(n7277), .B1(n532), .B2(n5824), .C1(n788), 
        .C2(n7278), .ZN(n7387) );
  AOI221_X1 U6495 ( .B1(n7279), .B2(n8167), .C1(n7280), .C2(n8103), .A(n7388), 
        .ZN(n7383) );
  OAI222_X1 U6496 ( .A1(n5039), .A2(n7282), .B1(n980), .B2(n5825), .C1(n5442), 
        .C2(n5816), .ZN(n7388) );
  AOI221_X1 U6497 ( .B1(n5833), .B2(DATAIN[13]), .C1(n7283), .C2(OUT2[13]), 
        .A(n7389), .ZN(n7382) );
  OAI22_X1 U6498 ( .A1(n4844), .A2(n5827), .B1(n5378), .B2(n7285), .ZN(n7389)
         );
  NAND4_X1 U6499 ( .A1(n7390), .A2(n7391), .A3(n7392), .A4(n7393), .ZN(n3650)
         );
  AOI221_X1 U6500 ( .B1(n7271), .B2(n5250), .C1(n7272), .C2(n4975), .A(n7394), 
        .ZN(n7393) );
  OAI222_X1 U6501 ( .A1(n1107), .A2(n5820), .B1(n1043), .B2(n5823), .C1(n1171), 
        .C2(n5815), .ZN(n7394) );
  AOI221_X1 U6502 ( .B1(n7274), .B2(n5315), .C1(n7275), .C2(n5104), .A(n7395), 
        .ZN(n7392) );
  OAI222_X1 U6503 ( .A1(n595), .A2(n7277), .B1(n531), .B2(n5824), .C1(n787), 
        .C2(n7278), .ZN(n7395) );
  AOI221_X1 U6504 ( .B1(n7279), .B2(n8166), .C1(n7280), .C2(n8102), .A(n7396), 
        .ZN(n7391) );
  OAI222_X1 U6505 ( .A1(n5040), .A2(n7282), .B1(n979), .B2(n5825), .C1(n5443), 
        .C2(n5816), .ZN(n7396) );
  AOI221_X1 U6506 ( .B1(n5833), .B2(DATAIN[14]), .C1(n7283), .C2(OUT2[14]), 
        .A(n7397), .ZN(n7390) );
  OAI22_X1 U6507 ( .A1(n4845), .A2(n5827), .B1(n5379), .B2(n7285), .ZN(n7397)
         );
  NAND4_X1 U6508 ( .A1(n7398), .A2(n7399), .A3(n7400), .A4(n7401), .ZN(n3649)
         );
  AOI221_X1 U6509 ( .B1(n7271), .B2(n5251), .C1(n7272), .C2(n4976), .A(n7402), 
        .ZN(n7401) );
  OAI222_X1 U6510 ( .A1(n1106), .A2(n5820), .B1(n1042), .B2(n5823), .C1(n1170), 
        .C2(n5815), .ZN(n7402) );
  AOI221_X1 U6511 ( .B1(n7274), .B2(n5316), .C1(n7275), .C2(n5105), .A(n7403), 
        .ZN(n7400) );
  OAI222_X1 U6512 ( .A1(n594), .A2(n7277), .B1(n530), .B2(n5824), .C1(n786), 
        .C2(n7278), .ZN(n7403) );
  AOI221_X1 U6513 ( .B1(n7279), .B2(n8165), .C1(n7280), .C2(n8101), .A(n7404), 
        .ZN(n7399) );
  OAI222_X1 U6514 ( .A1(n5041), .A2(n7282), .B1(n978), .B2(n5825), .C1(n5444), 
        .C2(n5816), .ZN(n7404) );
  AOI221_X1 U6515 ( .B1(n5833), .B2(DATAIN[15]), .C1(n7283), .C2(OUT2[15]), 
        .A(n7405), .ZN(n7398) );
  OAI22_X1 U6516 ( .A1(n4846), .A2(n5827), .B1(n5380), .B2(n7285), .ZN(n7405)
         );
  NAND4_X1 U6517 ( .A1(n7406), .A2(n7407), .A3(n7408), .A4(n7409), .ZN(n3648)
         );
  AOI221_X1 U6518 ( .B1(n7271), .B2(n5252), .C1(n7272), .C2(n4977), .A(n7410), 
        .ZN(n7409) );
  OAI222_X1 U6519 ( .A1(n1105), .A2(n5820), .B1(n1041), .B2(n5823), .C1(n1169), 
        .C2(n5815), .ZN(n7410) );
  AOI221_X1 U6520 ( .B1(n7274), .B2(n5317), .C1(n7275), .C2(n5106), .A(n7411), 
        .ZN(n7408) );
  OAI222_X1 U6521 ( .A1(n593), .A2(n7277), .B1(n529), .B2(n5824), .C1(n785), 
        .C2(n7278), .ZN(n7411) );
  AOI221_X1 U6522 ( .B1(n7279), .B2(n8164), .C1(n7280), .C2(n8100), .A(n7412), 
        .ZN(n7407) );
  OAI222_X1 U6523 ( .A1(n5042), .A2(n7282), .B1(n977), .B2(n5825), .C1(n5445), 
        .C2(n5816), .ZN(n7412) );
  AOI221_X1 U6524 ( .B1(n5833), .B2(DATAIN[16]), .C1(n7283), .C2(OUT2[16]), 
        .A(n7413), .ZN(n7406) );
  OAI22_X1 U6525 ( .A1(n4847), .A2(n5827), .B1(n5381), .B2(n7285), .ZN(n7413)
         );
  NAND4_X1 U6526 ( .A1(n7414), .A2(n7415), .A3(n7416), .A4(n7417), .ZN(n3647)
         );
  AOI221_X1 U6527 ( .B1(n7271), .B2(n5253), .C1(n7272), .C2(n4978), .A(n7418), 
        .ZN(n7417) );
  OAI222_X1 U6528 ( .A1(n1104), .A2(n5820), .B1(n1040), .B2(n5823), .C1(n1168), 
        .C2(n5815), .ZN(n7418) );
  AOI221_X1 U6529 ( .B1(n7274), .B2(n5318), .C1(n7275), .C2(n5107), .A(n7419), 
        .ZN(n7416) );
  OAI222_X1 U6530 ( .A1(n592), .A2(n7277), .B1(n528), .B2(n5824), .C1(n784), 
        .C2(n7278), .ZN(n7419) );
  AOI221_X1 U6531 ( .B1(n7279), .B2(n8163), .C1(n7280), .C2(n8099), .A(n7420), 
        .ZN(n7415) );
  OAI222_X1 U6532 ( .A1(n5043), .A2(n7282), .B1(n976), .B2(n5825), .C1(n5446), 
        .C2(n5816), .ZN(n7420) );
  AOI221_X1 U6533 ( .B1(n5833), .B2(DATAIN[17]), .C1(n7283), .C2(OUT2[17]), 
        .A(n7421), .ZN(n7414) );
  OAI22_X1 U6534 ( .A1(n4848), .A2(n5827), .B1(n5382), .B2(n7285), .ZN(n7421)
         );
  NAND4_X1 U6535 ( .A1(n7422), .A2(n7423), .A3(n7424), .A4(n7425), .ZN(n3646)
         );
  AOI221_X1 U6536 ( .B1(n7271), .B2(n5254), .C1(n7272), .C2(n4979), .A(n7426), 
        .ZN(n7425) );
  OAI222_X1 U6537 ( .A1(n1103), .A2(n5820), .B1(n1039), .B2(n5823), .C1(n1167), 
        .C2(n5815), .ZN(n7426) );
  AOI221_X1 U6538 ( .B1(n7274), .B2(n5319), .C1(n7275), .C2(n5108), .A(n7427), 
        .ZN(n7424) );
  OAI222_X1 U6539 ( .A1(n591), .A2(n7277), .B1(n527), .B2(n5824), .C1(n783), 
        .C2(n7278), .ZN(n7427) );
  AOI221_X1 U6540 ( .B1(n7279), .B2(n8162), .C1(n7280), .C2(n8098), .A(n7428), 
        .ZN(n7423) );
  OAI222_X1 U6541 ( .A1(n5044), .A2(n7282), .B1(n975), .B2(n5825), .C1(n5447), 
        .C2(n5816), .ZN(n7428) );
  AOI221_X1 U6542 ( .B1(n5833), .B2(DATAIN[18]), .C1(n7283), .C2(OUT2[18]), 
        .A(n7429), .ZN(n7422) );
  OAI22_X1 U6543 ( .A1(n4849), .A2(n5827), .B1(n5383), .B2(n7285), .ZN(n7429)
         );
  NAND4_X1 U6544 ( .A1(n7430), .A2(n7431), .A3(n7432), .A4(n7433), .ZN(n3645)
         );
  AOI221_X1 U6545 ( .B1(n7271), .B2(n5255), .C1(n7272), .C2(n4980), .A(n7434), 
        .ZN(n7433) );
  OAI222_X1 U6546 ( .A1(n1102), .A2(n5820), .B1(n1038), .B2(n5823), .C1(n1166), 
        .C2(n5815), .ZN(n7434) );
  AOI221_X1 U6547 ( .B1(n7274), .B2(n5320), .C1(n7275), .C2(n5109), .A(n7435), 
        .ZN(n7432) );
  OAI222_X1 U6548 ( .A1(n590), .A2(n7277), .B1(n526), .B2(n5824), .C1(n782), 
        .C2(n7278), .ZN(n7435) );
  AOI221_X1 U6549 ( .B1(n7279), .B2(n8161), .C1(n7280), .C2(n8097), .A(n7436), 
        .ZN(n7431) );
  OAI222_X1 U6550 ( .A1(n5045), .A2(n7282), .B1(n974), .B2(n5825), .C1(n5448), 
        .C2(n5816), .ZN(n7436) );
  AOI221_X1 U6551 ( .B1(n5833), .B2(DATAIN[19]), .C1(n7283), .C2(OUT2[19]), 
        .A(n7437), .ZN(n7430) );
  OAI22_X1 U6552 ( .A1(n4850), .A2(n5827), .B1(n5384), .B2(n7285), .ZN(n7437)
         );
  NAND4_X1 U6553 ( .A1(n7438), .A2(n7439), .A3(n7440), .A4(n7441), .ZN(n3644)
         );
  AOI221_X1 U6554 ( .B1(n7271), .B2(n5256), .C1(n7272), .C2(n4981), .A(n7442), 
        .ZN(n7441) );
  OAI222_X1 U6555 ( .A1(n1101), .A2(n5820), .B1(n1037), .B2(n5823), .C1(n1165), 
        .C2(n5815), .ZN(n7442) );
  AOI221_X1 U6556 ( .B1(n7274), .B2(n5321), .C1(n7275), .C2(n5110), .A(n7443), 
        .ZN(n7440) );
  OAI222_X1 U6557 ( .A1(n589), .A2(n7277), .B1(n525), .B2(n5824), .C1(n781), 
        .C2(n7278), .ZN(n7443) );
  AOI221_X1 U6558 ( .B1(n7279), .B2(n8160), .C1(n7280), .C2(n8096), .A(n7444), 
        .ZN(n7439) );
  OAI222_X1 U6559 ( .A1(n5046), .A2(n7282), .B1(n973), .B2(n5825), .C1(n5449), 
        .C2(n5816), .ZN(n7444) );
  AOI221_X1 U6560 ( .B1(n5833), .B2(DATAIN[20]), .C1(n7283), .C2(OUT2[20]), 
        .A(n7445), .ZN(n7438) );
  OAI22_X1 U6561 ( .A1(n4851), .A2(n5827), .B1(n5385), .B2(n7285), .ZN(n7445)
         );
  NAND4_X1 U6562 ( .A1(n7446), .A2(n7447), .A3(n7448), .A4(n7449), .ZN(n3643)
         );
  AOI221_X1 U6563 ( .B1(n7271), .B2(n5257), .C1(n7272), .C2(n4982), .A(n7450), 
        .ZN(n7449) );
  OAI222_X1 U6564 ( .A1(n1100), .A2(n5820), .B1(n1036), .B2(n5823), .C1(n1164), 
        .C2(n5815), .ZN(n7450) );
  AOI221_X1 U6565 ( .B1(n7274), .B2(n5322), .C1(n7275), .C2(n5111), .A(n7451), 
        .ZN(n7448) );
  OAI222_X1 U6566 ( .A1(n588), .A2(n7277), .B1(n524), .B2(n5824), .C1(n780), 
        .C2(n7278), .ZN(n7451) );
  AOI221_X1 U6567 ( .B1(n7279), .B2(n8159), .C1(n7280), .C2(n8095), .A(n7452), 
        .ZN(n7447) );
  OAI222_X1 U6568 ( .A1(n5047), .A2(n7282), .B1(n972), .B2(n5825), .C1(n5450), 
        .C2(n5816), .ZN(n7452) );
  AOI221_X1 U6569 ( .B1(n5833), .B2(DATAIN[21]), .C1(n7283), .C2(OUT2[21]), 
        .A(n7453), .ZN(n7446) );
  OAI22_X1 U6570 ( .A1(n4852), .A2(n5827), .B1(n5386), .B2(n7285), .ZN(n7453)
         );
  NAND4_X1 U6571 ( .A1(n7454), .A2(n7455), .A3(n7456), .A4(n7457), .ZN(n3642)
         );
  AOI221_X1 U6572 ( .B1(n7271), .B2(n5258), .C1(n7272), .C2(n4983), .A(n7458), 
        .ZN(n7457) );
  OAI222_X1 U6573 ( .A1(n1099), .A2(n5820), .B1(n1035), .B2(n5823), .C1(n1163), 
        .C2(n5815), .ZN(n7458) );
  AOI221_X1 U6574 ( .B1(n7274), .B2(n5323), .C1(n7275), .C2(n5112), .A(n7459), 
        .ZN(n7456) );
  OAI222_X1 U6575 ( .A1(n587), .A2(n7277), .B1(n523), .B2(n5824), .C1(n779), 
        .C2(n7278), .ZN(n7459) );
  AOI221_X1 U6576 ( .B1(n7279), .B2(n8158), .C1(n7280), .C2(n8094), .A(n7460), 
        .ZN(n7455) );
  OAI222_X1 U6577 ( .A1(n5048), .A2(n7282), .B1(n971), .B2(n5825), .C1(n5451), 
        .C2(n5816), .ZN(n7460) );
  AOI221_X1 U6578 ( .B1(n5833), .B2(DATAIN[22]), .C1(n7283), .C2(OUT2[22]), 
        .A(n7461), .ZN(n7454) );
  OAI22_X1 U6579 ( .A1(n4853), .A2(n5827), .B1(n5387), .B2(n7285), .ZN(n7461)
         );
  NAND4_X1 U6580 ( .A1(n7462), .A2(n7463), .A3(n7464), .A4(n7465), .ZN(n3641)
         );
  AOI221_X1 U6581 ( .B1(n7271), .B2(n5259), .C1(n7272), .C2(n4984), .A(n7466), 
        .ZN(n7465) );
  OAI222_X1 U6582 ( .A1(n1098), .A2(n5820), .B1(n1034), .B2(n5823), .C1(n1162), 
        .C2(n5815), .ZN(n7466) );
  AOI221_X1 U6583 ( .B1(n7274), .B2(n5324), .C1(n7275), .C2(n5113), .A(n7467), 
        .ZN(n7464) );
  OAI222_X1 U6584 ( .A1(n586), .A2(n7277), .B1(n522), .B2(n5824), .C1(n778), 
        .C2(n7278), .ZN(n7467) );
  AOI221_X1 U6585 ( .B1(n7279), .B2(n8157), .C1(n7280), .C2(n8093), .A(n7468), 
        .ZN(n7463) );
  OAI222_X1 U6586 ( .A1(n5049), .A2(n7282), .B1(n970), .B2(n5825), .C1(n5452), 
        .C2(n5816), .ZN(n7468) );
  AOI221_X1 U6587 ( .B1(n5833), .B2(DATAIN[23]), .C1(n7283), .C2(OUT2[23]), 
        .A(n7469), .ZN(n7462) );
  OAI22_X1 U6588 ( .A1(n4854), .A2(n5827), .B1(n5388), .B2(n7285), .ZN(n7469)
         );
  NAND4_X1 U6589 ( .A1(n7470), .A2(n7471), .A3(n7472), .A4(n7473), .ZN(n3640)
         );
  AOI221_X1 U6590 ( .B1(n7271), .B2(n5260), .C1(n7272), .C2(n4985), .A(n7474), 
        .ZN(n7473) );
  OAI222_X1 U6591 ( .A1(n1097), .A2(n5820), .B1(n1033), .B2(n5823), .C1(n1161), 
        .C2(n5815), .ZN(n7474) );
  AOI221_X1 U6592 ( .B1(n7274), .B2(n5325), .C1(n7275), .C2(n5114), .A(n7475), 
        .ZN(n7472) );
  OAI222_X1 U6593 ( .A1(n585), .A2(n7277), .B1(n521), .B2(n5824), .C1(n777), 
        .C2(n7278), .ZN(n7475) );
  AOI221_X1 U6594 ( .B1(n7279), .B2(n8156), .C1(n7280), .C2(n8092), .A(n7476), 
        .ZN(n7471) );
  OAI222_X1 U6595 ( .A1(n5050), .A2(n7282), .B1(n969), .B2(n5825), .C1(n5453), 
        .C2(n5816), .ZN(n7476) );
  AOI221_X1 U6596 ( .B1(n5833), .B2(DATAIN[24]), .C1(n7283), .C2(OUT2[24]), 
        .A(n7477), .ZN(n7470) );
  OAI22_X1 U6597 ( .A1(n4855), .A2(n5827), .B1(n5389), .B2(n7285), .ZN(n7477)
         );
  NAND4_X1 U6598 ( .A1(n7478), .A2(n7479), .A3(n7480), .A4(n7481), .ZN(n3639)
         );
  AOI221_X1 U6599 ( .B1(n7271), .B2(n5261), .C1(n7272), .C2(n4986), .A(n7482), 
        .ZN(n7481) );
  OAI222_X1 U6600 ( .A1(n1096), .A2(n5820), .B1(n1032), .B2(n5823), .C1(n1160), 
        .C2(n5815), .ZN(n7482) );
  AOI221_X1 U6601 ( .B1(n7274), .B2(n5326), .C1(n7275), .C2(n5115), .A(n7483), 
        .ZN(n7480) );
  OAI222_X1 U6602 ( .A1(n584), .A2(n7277), .B1(n520), .B2(n5824), .C1(n776), 
        .C2(n7278), .ZN(n7483) );
  AOI221_X1 U6603 ( .B1(n7279), .B2(n8155), .C1(n7280), .C2(n8091), .A(n7484), 
        .ZN(n7479) );
  OAI222_X1 U6604 ( .A1(n5051), .A2(n7282), .B1(n968), .B2(n5825), .C1(n5454), 
        .C2(n5816), .ZN(n7484) );
  AOI221_X1 U6605 ( .B1(n5833), .B2(DATAIN[25]), .C1(n7283), .C2(OUT2[25]), 
        .A(n7485), .ZN(n7478) );
  OAI22_X1 U6606 ( .A1(n4856), .A2(n5827), .B1(n5390), .B2(n7285), .ZN(n7485)
         );
  NAND4_X1 U6607 ( .A1(n7486), .A2(n7487), .A3(n7488), .A4(n7489), .ZN(n3638)
         );
  AOI221_X1 U6608 ( .B1(n7271), .B2(n5262), .C1(n7272), .C2(n4987), .A(n7490), 
        .ZN(n7489) );
  OAI222_X1 U6609 ( .A1(n1095), .A2(n5820), .B1(n1031), .B2(n5823), .C1(n1159), 
        .C2(n5815), .ZN(n7490) );
  AOI221_X1 U6610 ( .B1(n7274), .B2(n5327), .C1(n7275), .C2(n5116), .A(n7491), 
        .ZN(n7488) );
  OAI222_X1 U6611 ( .A1(n583), .A2(n7277), .B1(n519), .B2(n5824), .C1(n775), 
        .C2(n7278), .ZN(n7491) );
  AOI221_X1 U6612 ( .B1(n7279), .B2(n8154), .C1(n7280), .C2(n8090), .A(n7492), 
        .ZN(n7487) );
  OAI222_X1 U6613 ( .A1(n5052), .A2(n7282), .B1(n967), .B2(n5825), .C1(n5455), 
        .C2(n5816), .ZN(n7492) );
  AOI221_X1 U6614 ( .B1(n5833), .B2(DATAIN[26]), .C1(n7283), .C2(OUT2[26]), 
        .A(n7493), .ZN(n7486) );
  OAI22_X1 U6615 ( .A1(n4857), .A2(n5827), .B1(n5391), .B2(n7285), .ZN(n7493)
         );
  NAND4_X1 U6616 ( .A1(n7494), .A2(n7495), .A3(n7496), .A4(n7497), .ZN(n3637)
         );
  AOI221_X1 U6617 ( .B1(n7271), .B2(n5263), .C1(n7272), .C2(n4988), .A(n7498), 
        .ZN(n7497) );
  OAI222_X1 U6618 ( .A1(n1094), .A2(n5820), .B1(n1030), .B2(n5823), .C1(n1158), 
        .C2(n5815), .ZN(n7498) );
  AOI221_X1 U6619 ( .B1(n7274), .B2(n5328), .C1(n7275), .C2(n5117), .A(n7499), 
        .ZN(n7496) );
  OAI222_X1 U6620 ( .A1(n582), .A2(n7277), .B1(n518), .B2(n5824), .C1(n774), 
        .C2(n7278), .ZN(n7499) );
  AOI221_X1 U6621 ( .B1(n7279), .B2(n8153), .C1(n7280), .C2(n8089), .A(n7500), 
        .ZN(n7495) );
  OAI222_X1 U6622 ( .A1(n5053), .A2(n7282), .B1(n966), .B2(n5825), .C1(n5456), 
        .C2(n5816), .ZN(n7500) );
  AOI221_X1 U6623 ( .B1(n5833), .B2(DATAIN[27]), .C1(n7283), .C2(OUT2[27]), 
        .A(n7501), .ZN(n7494) );
  OAI22_X1 U6624 ( .A1(n4858), .A2(n5827), .B1(n5392), .B2(n7285), .ZN(n7501)
         );
  NAND4_X1 U6625 ( .A1(n7502), .A2(n7503), .A3(n7504), .A4(n7505), .ZN(n3636)
         );
  AOI221_X1 U6626 ( .B1(n7271), .B2(n5264), .C1(n7272), .C2(n4989), .A(n7506), 
        .ZN(n7505) );
  OAI222_X1 U6627 ( .A1(n1093), .A2(n5820), .B1(n1029), .B2(n5823), .C1(n1157), 
        .C2(n5815), .ZN(n7506) );
  AOI221_X1 U6628 ( .B1(n7274), .B2(n5329), .C1(n7275), .C2(n5118), .A(n7507), 
        .ZN(n7504) );
  OAI222_X1 U6629 ( .A1(n581), .A2(n7277), .B1(n517), .B2(n5824), .C1(n773), 
        .C2(n7278), .ZN(n7507) );
  AOI221_X1 U6630 ( .B1(n7279), .B2(n8152), .C1(n7280), .C2(n8088), .A(n7508), 
        .ZN(n7503) );
  OAI222_X1 U6631 ( .A1(n5054), .A2(n7282), .B1(n965), .B2(n5825), .C1(n5457), 
        .C2(n5816), .ZN(n7508) );
  AOI221_X1 U6632 ( .B1(n5833), .B2(DATAIN[28]), .C1(n7283), .C2(OUT2[28]), 
        .A(n7509), .ZN(n7502) );
  OAI22_X1 U6633 ( .A1(n4859), .A2(n5827), .B1(n5393), .B2(n7285), .ZN(n7509)
         );
  NAND4_X1 U6634 ( .A1(n7510), .A2(n7511), .A3(n7512), .A4(n7513), .ZN(n3635)
         );
  AOI221_X1 U6635 ( .B1(n7271), .B2(n5265), .C1(n7272), .C2(n4990), .A(n7514), 
        .ZN(n7513) );
  OAI222_X1 U6636 ( .A1(n1092), .A2(n5820), .B1(n1028), .B2(n5823), .C1(n1156), 
        .C2(n5815), .ZN(n7514) );
  AOI221_X1 U6637 ( .B1(n7274), .B2(n5330), .C1(n7275), .C2(n5119), .A(n7515), 
        .ZN(n7512) );
  OAI222_X1 U6638 ( .A1(n580), .A2(n7277), .B1(n516), .B2(n5824), .C1(n772), 
        .C2(n7278), .ZN(n7515) );
  AOI221_X1 U6639 ( .B1(n7279), .B2(n8151), .C1(n7280), .C2(n8087), .A(n7516), 
        .ZN(n7511) );
  OAI222_X1 U6640 ( .A1(n5055), .A2(n7282), .B1(n964), .B2(n5825), .C1(n5458), 
        .C2(n5816), .ZN(n7516) );
  AOI221_X1 U6641 ( .B1(n5833), .B2(DATAIN[29]), .C1(n7283), .C2(OUT2[29]), 
        .A(n7517), .ZN(n7510) );
  OAI22_X1 U6642 ( .A1(n4860), .A2(n5827), .B1(n5394), .B2(n7285), .ZN(n7517)
         );
  NAND4_X1 U6643 ( .A1(n7518), .A2(n7519), .A3(n7520), .A4(n7521), .ZN(n3634)
         );
  AOI221_X1 U6644 ( .B1(n7271), .B2(n5266), .C1(n7272), .C2(n4991), .A(n7522), 
        .ZN(n7521) );
  OAI222_X1 U6645 ( .A1(n1091), .A2(n5820), .B1(n1027), .B2(n5823), .C1(n1155), 
        .C2(n5815), .ZN(n7522) );
  AOI221_X1 U6646 ( .B1(n7274), .B2(n5331), .C1(n7275), .C2(n5120), .A(n7523), 
        .ZN(n7520) );
  OAI222_X1 U6647 ( .A1(n579), .A2(n7277), .B1(n515), .B2(n5824), .C1(n771), 
        .C2(n7278), .ZN(n7523) );
  AOI221_X1 U6648 ( .B1(n7279), .B2(n8150), .C1(n7280), .C2(n8086), .A(n7524), 
        .ZN(n7519) );
  OAI222_X1 U6649 ( .A1(n5056), .A2(n7282), .B1(n963), .B2(n5825), .C1(n5459), 
        .C2(n5816), .ZN(n7524) );
  AOI221_X1 U6650 ( .B1(n5833), .B2(DATAIN[30]), .C1(n7283), .C2(OUT2[30]), 
        .A(n7525), .ZN(n7518) );
  OAI22_X1 U6651 ( .A1(n4861), .A2(n5827), .B1(n5395), .B2(n7285), .ZN(n7525)
         );
  NAND4_X1 U6652 ( .A1(n7526), .A2(n7527), .A3(n7528), .A4(n7529), .ZN(n3633)
         );
  AOI221_X1 U6653 ( .B1(n7271), .B2(n5267), .C1(n7272), .C2(n4992), .A(n7530), 
        .ZN(n7529) );
  OAI222_X1 U6654 ( .A1(n1090), .A2(n5820), .B1(n1026), .B2(n5823), .C1(n1154), 
        .C2(n5815), .ZN(n7530) );
  AOI221_X1 U6655 ( .B1(n7274), .B2(n5332), .C1(n7275), .C2(n5121), .A(n7531), 
        .ZN(n7528) );
  OAI222_X1 U6656 ( .A1(n578), .A2(n7277), .B1(n514), .B2(n5824), .C1(n770), 
        .C2(n7278), .ZN(n7531) );
  AOI221_X1 U6657 ( .B1(n7279), .B2(n8149), .C1(n7280), .C2(n8085), .A(n7532), 
        .ZN(n7527) );
  OAI222_X1 U6658 ( .A1(n5057), .A2(n7282), .B1(n962), .B2(n5825), .C1(n5460), 
        .C2(n5816), .ZN(n7532) );
  AOI221_X1 U6659 ( .B1(n5833), .B2(DATAIN[31]), .C1(n7283), .C2(OUT2[31]), 
        .A(n7533), .ZN(n7526) );
  OAI22_X1 U6660 ( .A1(n4862), .A2(n5827), .B1(n5396), .B2(n7285), .ZN(n7533)
         );
  NAND4_X1 U6661 ( .A1(n7534), .A2(n7535), .A3(n7536), .A4(n7537), .ZN(n3632)
         );
  AOI221_X1 U6662 ( .B1(n7271), .B2(n5268), .C1(n7272), .C2(n4993), .A(n7538), 
        .ZN(n7537) );
  OAI222_X1 U6663 ( .A1(n1089), .A2(n5820), .B1(n1025), .B2(n5823), .C1(n1153), 
        .C2(n5815), .ZN(n7538) );
  AOI221_X1 U6664 ( .B1(n7274), .B2(n5333), .C1(n7275), .C2(n5122), .A(n7539), 
        .ZN(n7536) );
  OAI222_X1 U6665 ( .A1(n577), .A2(n7277), .B1(n513), .B2(n5824), .C1(n769), 
        .C2(n7278), .ZN(n7539) );
  AOI221_X1 U6666 ( .B1(n7279), .B2(n8148), .C1(n7280), .C2(n8084), .A(n7540), 
        .ZN(n7535) );
  OAI222_X1 U6667 ( .A1(n5058), .A2(n7282), .B1(n961), .B2(n5825), .C1(n5461), 
        .C2(n5816), .ZN(n7540) );
  AOI221_X1 U6668 ( .B1(n5833), .B2(DATAIN[32]), .C1(n7283), .C2(OUT2[32]), 
        .A(n7541), .ZN(n7534) );
  OAI22_X1 U6669 ( .A1(n4863), .A2(n5827), .B1(n5397), .B2(n7285), .ZN(n7541)
         );
  NAND4_X1 U6670 ( .A1(n7542), .A2(n7543), .A3(n7544), .A4(n7545), .ZN(n3631)
         );
  AOI221_X1 U6671 ( .B1(n7271), .B2(n5269), .C1(n7272), .C2(n4994), .A(n7546), 
        .ZN(n7545) );
  OAI222_X1 U6672 ( .A1(n1088), .A2(n5820), .B1(n1024), .B2(n5823), .C1(n1152), 
        .C2(n5815), .ZN(n7546) );
  AOI221_X1 U6673 ( .B1(n7274), .B2(n5334), .C1(n7275), .C2(n5123), .A(n7547), 
        .ZN(n7544) );
  OAI222_X1 U6674 ( .A1(n576), .A2(n7277), .B1(n512), .B2(n5824), .C1(n768), 
        .C2(n7278), .ZN(n7547) );
  AOI221_X1 U6675 ( .B1(n7279), .B2(n8147), .C1(n7280), .C2(n8083), .A(n7548), 
        .ZN(n7543) );
  OAI222_X1 U6676 ( .A1(n5059), .A2(n7282), .B1(n960), .B2(n5825), .C1(n5462), 
        .C2(n5816), .ZN(n7548) );
  AOI221_X1 U6677 ( .B1(n5833), .B2(DATAIN[33]), .C1(n7283), .C2(OUT2[33]), 
        .A(n7549), .ZN(n7542) );
  OAI22_X1 U6678 ( .A1(n4864), .A2(n5827), .B1(n5398), .B2(n7285), .ZN(n7549)
         );
  NAND4_X1 U6679 ( .A1(n7550), .A2(n7551), .A3(n7552), .A4(n7553), .ZN(n3630)
         );
  AOI221_X1 U6680 ( .B1(n7271), .B2(n5270), .C1(n7272), .C2(n4995), .A(n7554), 
        .ZN(n7553) );
  OAI222_X1 U6681 ( .A1(n1087), .A2(n5820), .B1(n1023), .B2(n5823), .C1(n1151), 
        .C2(n5815), .ZN(n7554) );
  AOI221_X1 U6682 ( .B1(n7274), .B2(n5335), .C1(n7275), .C2(n5124), .A(n7555), 
        .ZN(n7552) );
  OAI222_X1 U6683 ( .A1(n575), .A2(n7277), .B1(n511), .B2(n5824), .C1(n767), 
        .C2(n7278), .ZN(n7555) );
  AOI221_X1 U6684 ( .B1(n7279), .B2(n8146), .C1(n7280), .C2(n8082), .A(n7556), 
        .ZN(n7551) );
  OAI222_X1 U6685 ( .A1(n5060), .A2(n7282), .B1(n959), .B2(n5825), .C1(n5463), 
        .C2(n5816), .ZN(n7556) );
  AOI221_X1 U6686 ( .B1(n5833), .B2(DATAIN[34]), .C1(n7283), .C2(OUT2[34]), 
        .A(n7557), .ZN(n7550) );
  OAI22_X1 U6687 ( .A1(n4865), .A2(n5827), .B1(n5399), .B2(n7285), .ZN(n7557)
         );
  NAND4_X1 U6688 ( .A1(n7558), .A2(n7559), .A3(n7560), .A4(n7561), .ZN(n3629)
         );
  AOI221_X1 U6689 ( .B1(n7271), .B2(n5271), .C1(n7272), .C2(n4996), .A(n7562), 
        .ZN(n7561) );
  OAI222_X1 U6690 ( .A1(n1086), .A2(n5820), .B1(n1022), .B2(n5823), .C1(n1150), 
        .C2(n5815), .ZN(n7562) );
  AOI221_X1 U6691 ( .B1(n7274), .B2(n5336), .C1(n7275), .C2(n5125), .A(n7563), 
        .ZN(n7560) );
  OAI222_X1 U6692 ( .A1(n574), .A2(n7277), .B1(n510), .B2(n5824), .C1(n766), 
        .C2(n7278), .ZN(n7563) );
  AOI221_X1 U6693 ( .B1(n7279), .B2(n8145), .C1(n7280), .C2(n8081), .A(n7564), 
        .ZN(n7559) );
  OAI222_X1 U6694 ( .A1(n5061), .A2(n7282), .B1(n958), .B2(n5825), .C1(n5464), 
        .C2(n5816), .ZN(n7564) );
  AOI221_X1 U6695 ( .B1(n5833), .B2(DATAIN[35]), .C1(n7283), .C2(OUT2[35]), 
        .A(n7565), .ZN(n7558) );
  OAI22_X1 U6696 ( .A1(n4866), .A2(n5827), .B1(n5400), .B2(n7285), .ZN(n7565)
         );
  NAND4_X1 U6697 ( .A1(n7566), .A2(n7567), .A3(n7568), .A4(n7569), .ZN(n3628)
         );
  AOI221_X1 U6698 ( .B1(n7271), .B2(n5272), .C1(n7272), .C2(n4997), .A(n7570), 
        .ZN(n7569) );
  OAI222_X1 U6699 ( .A1(n1085), .A2(n5820), .B1(n1021), .B2(n5823), .C1(n1149), 
        .C2(n5815), .ZN(n7570) );
  AOI221_X1 U6700 ( .B1(n7274), .B2(n5337), .C1(n7275), .C2(n5126), .A(n7571), 
        .ZN(n7568) );
  OAI222_X1 U6701 ( .A1(n573), .A2(n7277), .B1(n509), .B2(n5824), .C1(n765), 
        .C2(n7278), .ZN(n7571) );
  AOI221_X1 U6702 ( .B1(n7279), .B2(n8144), .C1(n7280), .C2(n8080), .A(n7572), 
        .ZN(n7567) );
  OAI222_X1 U6703 ( .A1(n5062), .A2(n7282), .B1(n957), .B2(n5825), .C1(n5465), 
        .C2(n5816), .ZN(n7572) );
  AOI221_X1 U6704 ( .B1(n5833), .B2(DATAIN[36]), .C1(n7283), .C2(OUT2[36]), 
        .A(n7573), .ZN(n7566) );
  OAI22_X1 U6705 ( .A1(n4867), .A2(n5827), .B1(n5401), .B2(n7285), .ZN(n7573)
         );
  NAND4_X1 U6706 ( .A1(n7574), .A2(n7575), .A3(n7576), .A4(n7577), .ZN(n3627)
         );
  AOI221_X1 U6707 ( .B1(n7271), .B2(n5273), .C1(n7272), .C2(n4998), .A(n7578), 
        .ZN(n7577) );
  OAI222_X1 U6708 ( .A1(n1084), .A2(n5820), .B1(n1020), .B2(n5823), .C1(n1148), 
        .C2(n5815), .ZN(n7578) );
  AOI221_X1 U6709 ( .B1(n7274), .B2(n5338), .C1(n7275), .C2(n5127), .A(n7579), 
        .ZN(n7576) );
  OAI222_X1 U6710 ( .A1(n572), .A2(n7277), .B1(n508), .B2(n5824), .C1(n764), 
        .C2(n7278), .ZN(n7579) );
  AOI221_X1 U6711 ( .B1(n7279), .B2(n8143), .C1(n7280), .C2(n8079), .A(n7580), 
        .ZN(n7575) );
  OAI222_X1 U6712 ( .A1(n5063), .A2(n7282), .B1(n956), .B2(n5825), .C1(n5466), 
        .C2(n5816), .ZN(n7580) );
  AOI221_X1 U6713 ( .B1(n5833), .B2(DATAIN[37]), .C1(n7283), .C2(OUT2[37]), 
        .A(n7581), .ZN(n7574) );
  OAI22_X1 U6714 ( .A1(n4868), .A2(n5827), .B1(n5402), .B2(n7285), .ZN(n7581)
         );
  NAND4_X1 U6715 ( .A1(n7582), .A2(n7583), .A3(n7584), .A4(n7585), .ZN(n3626)
         );
  AOI221_X1 U6716 ( .B1(n7271), .B2(n5274), .C1(n7272), .C2(n4999), .A(n7586), 
        .ZN(n7585) );
  OAI222_X1 U6717 ( .A1(n1083), .A2(n5820), .B1(n1019), .B2(n5823), .C1(n1147), 
        .C2(n5815), .ZN(n7586) );
  AOI221_X1 U6718 ( .B1(n7274), .B2(n5339), .C1(n7275), .C2(n5128), .A(n7587), 
        .ZN(n7584) );
  OAI222_X1 U6719 ( .A1(n571), .A2(n7277), .B1(n507), .B2(n5824), .C1(n763), 
        .C2(n7278), .ZN(n7587) );
  AOI221_X1 U6720 ( .B1(n7279), .B2(n8142), .C1(n7280), .C2(n8078), .A(n7588), 
        .ZN(n7583) );
  OAI222_X1 U6721 ( .A1(n5064), .A2(n7282), .B1(n955), .B2(n5825), .C1(n5467), 
        .C2(n5816), .ZN(n7588) );
  AOI221_X1 U6722 ( .B1(n5833), .B2(DATAIN[38]), .C1(n7283), .C2(OUT2[38]), 
        .A(n7589), .ZN(n7582) );
  OAI22_X1 U6723 ( .A1(n4869), .A2(n5827), .B1(n5403), .B2(n7285), .ZN(n7589)
         );
  NAND4_X1 U6724 ( .A1(n7590), .A2(n7591), .A3(n7592), .A4(n7593), .ZN(n3625)
         );
  AOI221_X1 U6725 ( .B1(n7271), .B2(n5275), .C1(n7272), .C2(n5000), .A(n7594), 
        .ZN(n7593) );
  OAI222_X1 U6726 ( .A1(n1082), .A2(n5820), .B1(n1018), .B2(n5823), .C1(n1146), 
        .C2(n5815), .ZN(n7594) );
  AOI221_X1 U6727 ( .B1(n7274), .B2(n5340), .C1(n7275), .C2(n5129), .A(n7595), 
        .ZN(n7592) );
  OAI222_X1 U6728 ( .A1(n570), .A2(n7277), .B1(n506), .B2(n5824), .C1(n762), 
        .C2(n7278), .ZN(n7595) );
  AOI221_X1 U6729 ( .B1(n7279), .B2(n8141), .C1(n7280), .C2(n8077), .A(n7596), 
        .ZN(n7591) );
  OAI222_X1 U6730 ( .A1(n5065), .A2(n7282), .B1(n954), .B2(n5825), .C1(n5468), 
        .C2(n5816), .ZN(n7596) );
  AOI221_X1 U6731 ( .B1(n5833), .B2(DATAIN[39]), .C1(n7283), .C2(OUT2[39]), 
        .A(n7597), .ZN(n7590) );
  OAI22_X1 U6732 ( .A1(n4870), .A2(n5827), .B1(n5404), .B2(n7285), .ZN(n7597)
         );
  NAND4_X1 U6733 ( .A1(n7598), .A2(n7599), .A3(n7600), .A4(n7601), .ZN(n3624)
         );
  AOI221_X1 U6734 ( .B1(n7271), .B2(n5276), .C1(n7272), .C2(n5001), .A(n7602), 
        .ZN(n7601) );
  OAI222_X1 U6735 ( .A1(n1081), .A2(n5820), .B1(n1017), .B2(n5823), .C1(n1145), 
        .C2(n5815), .ZN(n7602) );
  AOI221_X1 U6736 ( .B1(n7274), .B2(n5341), .C1(n7275), .C2(n5130), .A(n7603), 
        .ZN(n7600) );
  OAI222_X1 U6737 ( .A1(n569), .A2(n7277), .B1(n505), .B2(n5824), .C1(n761), 
        .C2(n7278), .ZN(n7603) );
  AOI221_X1 U6738 ( .B1(n7279), .B2(n8140), .C1(n7280), .C2(n8076), .A(n7604), 
        .ZN(n7599) );
  OAI222_X1 U6739 ( .A1(n5066), .A2(n7282), .B1(n953), .B2(n5825), .C1(n5469), 
        .C2(n5816), .ZN(n7604) );
  AOI221_X1 U6740 ( .B1(n5833), .B2(DATAIN[40]), .C1(n7283), .C2(OUT2[40]), 
        .A(n7605), .ZN(n7598) );
  OAI22_X1 U6741 ( .A1(n4871), .A2(n5827), .B1(n5405), .B2(n7285), .ZN(n7605)
         );
  NAND4_X1 U6742 ( .A1(n7606), .A2(n7607), .A3(n7608), .A4(n7609), .ZN(n3623)
         );
  AOI221_X1 U6743 ( .B1(n7271), .B2(n5277), .C1(n7272), .C2(n5002), .A(n7610), 
        .ZN(n7609) );
  OAI222_X1 U6744 ( .A1(n1080), .A2(n5820), .B1(n1016), .B2(n5823), .C1(n1144), 
        .C2(n5815), .ZN(n7610) );
  AOI221_X1 U6745 ( .B1(n7274), .B2(n5342), .C1(n7275), .C2(n5131), .A(n7611), 
        .ZN(n7608) );
  OAI222_X1 U6746 ( .A1(n568), .A2(n7277), .B1(n504), .B2(n5824), .C1(n760), 
        .C2(n7278), .ZN(n7611) );
  AOI221_X1 U6747 ( .B1(n7279), .B2(n8139), .C1(n7280), .C2(n8075), .A(n7612), 
        .ZN(n7607) );
  OAI222_X1 U6748 ( .A1(n5067), .A2(n7282), .B1(n952), .B2(n5825), .C1(n5470), 
        .C2(n5816), .ZN(n7612) );
  AOI221_X1 U6749 ( .B1(n5833), .B2(DATAIN[41]), .C1(n7283), .C2(OUT2[41]), 
        .A(n7613), .ZN(n7606) );
  OAI22_X1 U6750 ( .A1(n4872), .A2(n5827), .B1(n5406), .B2(n7285), .ZN(n7613)
         );
  NAND4_X1 U6751 ( .A1(n7614), .A2(n7615), .A3(n7616), .A4(n7617), .ZN(n3622)
         );
  AOI221_X1 U6752 ( .B1(n7271), .B2(n5278), .C1(n7272), .C2(n5003), .A(n7618), 
        .ZN(n7617) );
  OAI222_X1 U6753 ( .A1(n1079), .A2(n5820), .B1(n1015), .B2(n5823), .C1(n1143), 
        .C2(n5815), .ZN(n7618) );
  AOI221_X1 U6754 ( .B1(n7274), .B2(n5343), .C1(n7275), .C2(n5132), .A(n7619), 
        .ZN(n7616) );
  OAI222_X1 U6755 ( .A1(n567), .A2(n7277), .B1(n503), .B2(n5824), .C1(n759), 
        .C2(n7278), .ZN(n7619) );
  AOI221_X1 U6756 ( .B1(n7279), .B2(n8138), .C1(n7280), .C2(n8074), .A(n7620), 
        .ZN(n7615) );
  OAI222_X1 U6757 ( .A1(n5068), .A2(n7282), .B1(n951), .B2(n5825), .C1(n5471), 
        .C2(n5816), .ZN(n7620) );
  AOI221_X1 U6758 ( .B1(n5833), .B2(DATAIN[42]), .C1(n7283), .C2(OUT2[42]), 
        .A(n7621), .ZN(n7614) );
  OAI22_X1 U6759 ( .A1(n4873), .A2(n5827), .B1(n5407), .B2(n7285), .ZN(n7621)
         );
  NAND4_X1 U6760 ( .A1(n7622), .A2(n7623), .A3(n7624), .A4(n7625), .ZN(n3621)
         );
  AOI221_X1 U6761 ( .B1(n7271), .B2(n5279), .C1(n7272), .C2(n5004), .A(n7626), 
        .ZN(n7625) );
  OAI222_X1 U6762 ( .A1(n1078), .A2(n5820), .B1(n1014), .B2(n5823), .C1(n1142), 
        .C2(n5815), .ZN(n7626) );
  AOI221_X1 U6763 ( .B1(n7274), .B2(n5344), .C1(n7275), .C2(n5133), .A(n7627), 
        .ZN(n7624) );
  OAI222_X1 U6764 ( .A1(n566), .A2(n7277), .B1(n502), .B2(n5824), .C1(n758), 
        .C2(n7278), .ZN(n7627) );
  AOI221_X1 U6765 ( .B1(n7279), .B2(n8137), .C1(n7280), .C2(n8073), .A(n7628), 
        .ZN(n7623) );
  OAI222_X1 U6766 ( .A1(n5069), .A2(n7282), .B1(n950), .B2(n5825), .C1(n5472), 
        .C2(n5816), .ZN(n7628) );
  AOI221_X1 U6767 ( .B1(n5833), .B2(DATAIN[43]), .C1(n7283), .C2(OUT2[43]), 
        .A(n7629), .ZN(n7622) );
  OAI22_X1 U6768 ( .A1(n4874), .A2(n5827), .B1(n5408), .B2(n7285), .ZN(n7629)
         );
  NAND4_X1 U6769 ( .A1(n7630), .A2(n7631), .A3(n7632), .A4(n7633), .ZN(n3620)
         );
  AOI221_X1 U6770 ( .B1(n7271), .B2(n5280), .C1(n7272), .C2(n5005), .A(n7634), 
        .ZN(n7633) );
  OAI222_X1 U6771 ( .A1(n1077), .A2(n5820), .B1(n1013), .B2(n5823), .C1(n1141), 
        .C2(n5815), .ZN(n7634) );
  AOI221_X1 U6772 ( .B1(n7274), .B2(n5345), .C1(n7275), .C2(n5134), .A(n7635), 
        .ZN(n7632) );
  OAI222_X1 U6773 ( .A1(n565), .A2(n7277), .B1(n501), .B2(n5824), .C1(n757), 
        .C2(n7278), .ZN(n7635) );
  AOI221_X1 U6774 ( .B1(n7279), .B2(n8136), .C1(n7280), .C2(n8072), .A(n7636), 
        .ZN(n7631) );
  OAI222_X1 U6775 ( .A1(n5070), .A2(n7282), .B1(n949), .B2(n5825), .C1(n5473), 
        .C2(n5816), .ZN(n7636) );
  AOI221_X1 U6776 ( .B1(n5833), .B2(DATAIN[44]), .C1(n7283), .C2(OUT2[44]), 
        .A(n7637), .ZN(n7630) );
  OAI22_X1 U6777 ( .A1(n4875), .A2(n5827), .B1(n5409), .B2(n7285), .ZN(n7637)
         );
  NAND4_X1 U6778 ( .A1(n7638), .A2(n7639), .A3(n7640), .A4(n7641), .ZN(n3619)
         );
  AOI221_X1 U6779 ( .B1(n7271), .B2(n5281), .C1(n7272), .C2(n5006), .A(n7642), 
        .ZN(n7641) );
  OAI222_X1 U6780 ( .A1(n1076), .A2(n5820), .B1(n1012), .B2(n5823), .C1(n1140), 
        .C2(n5815), .ZN(n7642) );
  AOI221_X1 U6781 ( .B1(n7274), .B2(n5346), .C1(n7275), .C2(n5135), .A(n7643), 
        .ZN(n7640) );
  OAI222_X1 U6782 ( .A1(n564), .A2(n7277), .B1(n500), .B2(n5824), .C1(n756), 
        .C2(n7278), .ZN(n7643) );
  AOI221_X1 U6783 ( .B1(n7279), .B2(n8135), .C1(n7280), .C2(n8071), .A(n7644), 
        .ZN(n7639) );
  OAI222_X1 U6784 ( .A1(n5071), .A2(n7282), .B1(n948), .B2(n5825), .C1(n5474), 
        .C2(n5816), .ZN(n7644) );
  AOI221_X1 U6785 ( .B1(n5833), .B2(DATAIN[45]), .C1(n7283), .C2(OUT2[45]), 
        .A(n7645), .ZN(n7638) );
  OAI22_X1 U6786 ( .A1(n4876), .A2(n5827), .B1(n5410), .B2(n7285), .ZN(n7645)
         );
  NAND4_X1 U6787 ( .A1(n7646), .A2(n7647), .A3(n7648), .A4(n7649), .ZN(n3618)
         );
  AOI221_X1 U6788 ( .B1(n7271), .B2(n5282), .C1(n7272), .C2(n5007), .A(n7650), 
        .ZN(n7649) );
  OAI222_X1 U6789 ( .A1(n1075), .A2(n5820), .B1(n1011), .B2(n5823), .C1(n1139), 
        .C2(n5815), .ZN(n7650) );
  AOI221_X1 U6790 ( .B1(n7274), .B2(n5347), .C1(n7275), .C2(n5136), .A(n7651), 
        .ZN(n7648) );
  OAI222_X1 U6791 ( .A1(n563), .A2(n7277), .B1(n499), .B2(n5824), .C1(n755), 
        .C2(n7278), .ZN(n7651) );
  AOI221_X1 U6792 ( .B1(n7279), .B2(n8134), .C1(n7280), .C2(n8070), .A(n7652), 
        .ZN(n7647) );
  OAI222_X1 U6793 ( .A1(n5072), .A2(n7282), .B1(n947), .B2(n5825), .C1(n5475), 
        .C2(n5816), .ZN(n7652) );
  AOI221_X1 U6794 ( .B1(n5833), .B2(DATAIN[46]), .C1(n7283), .C2(OUT2[46]), 
        .A(n7653), .ZN(n7646) );
  OAI22_X1 U6795 ( .A1(n4877), .A2(n5827), .B1(n5411), .B2(n7285), .ZN(n7653)
         );
  NAND4_X1 U6796 ( .A1(n7654), .A2(n7655), .A3(n7656), .A4(n7657), .ZN(n3617)
         );
  AOI221_X1 U6797 ( .B1(n7271), .B2(n5283), .C1(n7272), .C2(n5008), .A(n7658), 
        .ZN(n7657) );
  OAI222_X1 U6798 ( .A1(n1074), .A2(n5820), .B1(n1010), .B2(n5823), .C1(n1138), 
        .C2(n5815), .ZN(n7658) );
  AOI221_X1 U6799 ( .B1(n7274), .B2(n5348), .C1(n7275), .C2(n5137), .A(n7659), 
        .ZN(n7656) );
  OAI222_X1 U6800 ( .A1(n562), .A2(n7277), .B1(n498), .B2(n5824), .C1(n754), 
        .C2(n7278), .ZN(n7659) );
  AOI221_X1 U6801 ( .B1(n7279), .B2(n8133), .C1(n7280), .C2(n8069), .A(n7660), 
        .ZN(n7655) );
  OAI222_X1 U6802 ( .A1(n5073), .A2(n7282), .B1(n946), .B2(n5825), .C1(n5476), 
        .C2(n5816), .ZN(n7660) );
  AOI221_X1 U6803 ( .B1(n5833), .B2(DATAIN[47]), .C1(n7283), .C2(OUT2[47]), 
        .A(n7661), .ZN(n7654) );
  OAI22_X1 U6804 ( .A1(n4878), .A2(n5827), .B1(n5412), .B2(n7285), .ZN(n7661)
         );
  NAND4_X1 U6805 ( .A1(n7662), .A2(n7663), .A3(n7664), .A4(n7665), .ZN(n3616)
         );
  AOI221_X1 U6806 ( .B1(n7271), .B2(n5284), .C1(n7272), .C2(n5009), .A(n7666), 
        .ZN(n7665) );
  OAI222_X1 U6807 ( .A1(n1073), .A2(n5820), .B1(n1009), .B2(n5823), .C1(n1137), 
        .C2(n5815), .ZN(n7666) );
  AOI221_X1 U6808 ( .B1(n7274), .B2(n5349), .C1(n7275), .C2(n5138), .A(n7667), 
        .ZN(n7664) );
  OAI222_X1 U6809 ( .A1(n561), .A2(n7277), .B1(n497), .B2(n5824), .C1(n753), 
        .C2(n7278), .ZN(n7667) );
  AOI221_X1 U6810 ( .B1(n7279), .B2(n8132), .C1(n7280), .C2(n8068), .A(n7668), 
        .ZN(n7663) );
  OAI222_X1 U6811 ( .A1(n5074), .A2(n7282), .B1(n945), .B2(n5825), .C1(n5477), 
        .C2(n5816), .ZN(n7668) );
  AOI221_X1 U6812 ( .B1(n5833), .B2(DATAIN[48]), .C1(n7283), .C2(OUT2[48]), 
        .A(n7669), .ZN(n7662) );
  OAI22_X1 U6813 ( .A1(n4879), .A2(n5827), .B1(n5413), .B2(n7285), .ZN(n7669)
         );
  NAND4_X1 U6814 ( .A1(n7670), .A2(n7671), .A3(n7672), .A4(n7673), .ZN(n3615)
         );
  AOI221_X1 U6815 ( .B1(n7271), .B2(n5285), .C1(n7272), .C2(n5010), .A(n7674), 
        .ZN(n7673) );
  OAI222_X1 U6816 ( .A1(n1072), .A2(n5820), .B1(n1008), .B2(n5823), .C1(n1136), 
        .C2(n5815), .ZN(n7674) );
  AOI221_X1 U6817 ( .B1(n7274), .B2(n5350), .C1(n7275), .C2(n5139), .A(n7675), 
        .ZN(n7672) );
  OAI222_X1 U6818 ( .A1(n560), .A2(n7277), .B1(n496), .B2(n5824), .C1(n752), 
        .C2(n7278), .ZN(n7675) );
  AOI221_X1 U6819 ( .B1(n7279), .B2(n8131), .C1(n7280), .C2(n8067), .A(n7676), 
        .ZN(n7671) );
  OAI222_X1 U6820 ( .A1(n5075), .A2(n7282), .B1(n944), .B2(n5825), .C1(n5478), 
        .C2(n5816), .ZN(n7676) );
  AOI221_X1 U6821 ( .B1(n5833), .B2(DATAIN[49]), .C1(n7283), .C2(OUT2[49]), 
        .A(n7677), .ZN(n7670) );
  OAI22_X1 U6822 ( .A1(n4880), .A2(n5827), .B1(n5414), .B2(n7285), .ZN(n7677)
         );
  NAND4_X1 U6823 ( .A1(n7678), .A2(n7679), .A3(n7680), .A4(n7681), .ZN(n3614)
         );
  AOI221_X1 U6824 ( .B1(n7271), .B2(n5286), .C1(n7272), .C2(n5011), .A(n7682), 
        .ZN(n7681) );
  OAI222_X1 U6825 ( .A1(n1071), .A2(n5820), .B1(n1007), .B2(n5823), .C1(n1135), 
        .C2(n5815), .ZN(n7682) );
  AOI221_X1 U6826 ( .B1(n7274), .B2(n5351), .C1(n7275), .C2(n5140), .A(n7683), 
        .ZN(n7680) );
  OAI222_X1 U6827 ( .A1(n559), .A2(n7277), .B1(n495), .B2(n5824), .C1(n751), 
        .C2(n7278), .ZN(n7683) );
  AOI221_X1 U6828 ( .B1(n7279), .B2(n8130), .C1(n7280), .C2(n8066), .A(n7684), 
        .ZN(n7679) );
  OAI222_X1 U6829 ( .A1(n5076), .A2(n7282), .B1(n943), .B2(n5825), .C1(n5479), 
        .C2(n5816), .ZN(n7684) );
  AOI221_X1 U6830 ( .B1(n5833), .B2(DATAIN[50]), .C1(n7283), .C2(OUT2[50]), 
        .A(n7685), .ZN(n7678) );
  OAI22_X1 U6831 ( .A1(n4881), .A2(n5827), .B1(n5415), .B2(n7285), .ZN(n7685)
         );
  NAND4_X1 U6832 ( .A1(n7686), .A2(n7687), .A3(n7688), .A4(n7689), .ZN(n3613)
         );
  AOI221_X1 U6833 ( .B1(n7271), .B2(n5287), .C1(n7272), .C2(n5012), .A(n7690), 
        .ZN(n7689) );
  OAI222_X1 U6834 ( .A1(n1070), .A2(n5820), .B1(n1006), .B2(n5823), .C1(n1134), 
        .C2(n5815), .ZN(n7690) );
  AOI221_X1 U6835 ( .B1(n7274), .B2(n5352), .C1(n7275), .C2(n5141), .A(n7691), 
        .ZN(n7688) );
  OAI222_X1 U6836 ( .A1(n558), .A2(n7277), .B1(n494), .B2(n5824), .C1(n750), 
        .C2(n7278), .ZN(n7691) );
  AOI221_X1 U6837 ( .B1(n7279), .B2(n8129), .C1(n7280), .C2(n8065), .A(n7692), 
        .ZN(n7687) );
  OAI222_X1 U6838 ( .A1(n5077), .A2(n7282), .B1(n942), .B2(n5825), .C1(n5480), 
        .C2(n5816), .ZN(n7692) );
  AOI221_X1 U6839 ( .B1(n5833), .B2(DATAIN[51]), .C1(n7283), .C2(OUT2[51]), 
        .A(n7693), .ZN(n7686) );
  OAI22_X1 U6840 ( .A1(n4882), .A2(n5827), .B1(n5416), .B2(n7285), .ZN(n7693)
         );
  NAND4_X1 U6841 ( .A1(n7694), .A2(n7695), .A3(n7696), .A4(n7697), .ZN(n3612)
         );
  AOI221_X1 U6842 ( .B1(n7271), .B2(n5288), .C1(n7272), .C2(n5013), .A(n7698), 
        .ZN(n7697) );
  OAI222_X1 U6843 ( .A1(n1069), .A2(n5820), .B1(n1005), .B2(n5823), .C1(n1133), 
        .C2(n5815), .ZN(n7698) );
  AOI221_X1 U6844 ( .B1(n7274), .B2(n5353), .C1(n7275), .C2(n5142), .A(n7699), 
        .ZN(n7696) );
  OAI222_X1 U6845 ( .A1(n557), .A2(n7277), .B1(n493), .B2(n5824), .C1(n749), 
        .C2(n7278), .ZN(n7699) );
  AOI221_X1 U6846 ( .B1(n7279), .B2(n8128), .C1(n7280), .C2(n8064), .A(n7700), 
        .ZN(n7695) );
  OAI222_X1 U6847 ( .A1(n5078), .A2(n7282), .B1(n941), .B2(n5825), .C1(n5481), 
        .C2(n5816), .ZN(n7700) );
  AOI221_X1 U6848 ( .B1(n5833), .B2(DATAIN[52]), .C1(n7283), .C2(OUT2[52]), 
        .A(n7701), .ZN(n7694) );
  OAI22_X1 U6849 ( .A1(n4883), .A2(n5827), .B1(n5417), .B2(n7285), .ZN(n7701)
         );
  NAND4_X1 U6850 ( .A1(n7702), .A2(n7703), .A3(n7704), .A4(n7705), .ZN(n3611)
         );
  AOI221_X1 U6851 ( .B1(n7271), .B2(n5289), .C1(n7272), .C2(n5014), .A(n7706), 
        .ZN(n7705) );
  OAI222_X1 U6852 ( .A1(n1068), .A2(n5820), .B1(n1004), .B2(n5823), .C1(n1132), 
        .C2(n5815), .ZN(n7706) );
  AOI221_X1 U6853 ( .B1(n7274), .B2(n5354), .C1(n7275), .C2(n5143), .A(n7707), 
        .ZN(n7704) );
  OAI222_X1 U6854 ( .A1(n556), .A2(n7277), .B1(n492), .B2(n5824), .C1(n748), 
        .C2(n7278), .ZN(n7707) );
  AOI221_X1 U6855 ( .B1(n7279), .B2(n8127), .C1(n7280), .C2(n8063), .A(n7708), 
        .ZN(n7703) );
  OAI222_X1 U6856 ( .A1(n5079), .A2(n7282), .B1(n940), .B2(n5825), .C1(n5482), 
        .C2(n5816), .ZN(n7708) );
  AOI221_X1 U6857 ( .B1(n5833), .B2(DATAIN[53]), .C1(n7283), .C2(OUT2[53]), 
        .A(n7709), .ZN(n7702) );
  OAI22_X1 U6858 ( .A1(n4884), .A2(n5827), .B1(n5418), .B2(n7285), .ZN(n7709)
         );
  NAND4_X1 U6859 ( .A1(n7710), .A2(n7711), .A3(n7712), .A4(n7713), .ZN(n3610)
         );
  AOI221_X1 U6860 ( .B1(n7271), .B2(n5290), .C1(n7272), .C2(n5015), .A(n7714), 
        .ZN(n7713) );
  OAI222_X1 U6861 ( .A1(n1067), .A2(n5820), .B1(n1003), .B2(n5823), .C1(n1131), 
        .C2(n5815), .ZN(n7714) );
  AOI221_X1 U6862 ( .B1(n7274), .B2(n5355), .C1(n7275), .C2(n5144), .A(n7715), 
        .ZN(n7712) );
  OAI222_X1 U6863 ( .A1(n555), .A2(n7277), .B1(n491), .B2(n5824), .C1(n747), 
        .C2(n7278), .ZN(n7715) );
  AOI221_X1 U6864 ( .B1(n7279), .B2(n8126), .C1(n7280), .C2(n8062), .A(n7716), 
        .ZN(n7711) );
  OAI222_X1 U6865 ( .A1(n5080), .A2(n7282), .B1(n939), .B2(n5825), .C1(n5483), 
        .C2(n5816), .ZN(n7716) );
  AOI221_X1 U6866 ( .B1(n5833), .B2(DATAIN[54]), .C1(n7283), .C2(OUT2[54]), 
        .A(n7717), .ZN(n7710) );
  OAI22_X1 U6867 ( .A1(n4885), .A2(n5827), .B1(n5419), .B2(n7285), .ZN(n7717)
         );
  NAND4_X1 U6868 ( .A1(n7718), .A2(n7719), .A3(n7720), .A4(n7721), .ZN(n3609)
         );
  AOI221_X1 U6869 ( .B1(n7271), .B2(n5291), .C1(n7272), .C2(n5016), .A(n7722), 
        .ZN(n7721) );
  OAI222_X1 U6870 ( .A1(n1066), .A2(n5820), .B1(n1002), .B2(n5823), .C1(n1130), 
        .C2(n5815), .ZN(n7722) );
  AOI221_X1 U6871 ( .B1(n7274), .B2(n5356), .C1(n7275), .C2(n5145), .A(n7723), 
        .ZN(n7720) );
  OAI222_X1 U6872 ( .A1(n554), .A2(n7277), .B1(n490), .B2(n5824), .C1(n746), 
        .C2(n7278), .ZN(n7723) );
  AOI221_X1 U6873 ( .B1(n7279), .B2(n8125), .C1(n7280), .C2(n8061), .A(n7724), 
        .ZN(n7719) );
  OAI222_X1 U6874 ( .A1(n5081), .A2(n7282), .B1(n938), .B2(n5825), .C1(n5484), 
        .C2(n5816), .ZN(n7724) );
  AOI221_X1 U6875 ( .B1(n5833), .B2(DATAIN[55]), .C1(n7283), .C2(OUT2[55]), 
        .A(n7725), .ZN(n7718) );
  OAI22_X1 U6876 ( .A1(n4886), .A2(n5827), .B1(n5420), .B2(n7285), .ZN(n7725)
         );
  NAND4_X1 U6877 ( .A1(n7726), .A2(n7727), .A3(n7728), .A4(n7729), .ZN(n3608)
         );
  AOI221_X1 U6878 ( .B1(n7271), .B2(n5292), .C1(n7272), .C2(n5017), .A(n7730), 
        .ZN(n7729) );
  OAI222_X1 U6879 ( .A1(n1065), .A2(n5820), .B1(n1001), .B2(n5823), .C1(n1129), 
        .C2(n5815), .ZN(n7730) );
  AOI221_X1 U6880 ( .B1(n7274), .B2(n5357), .C1(n7275), .C2(n5146), .A(n7731), 
        .ZN(n7728) );
  OAI222_X1 U6881 ( .A1(n553), .A2(n7277), .B1(n489), .B2(n5824), .C1(n745), 
        .C2(n7278), .ZN(n7731) );
  AOI221_X1 U6882 ( .B1(n7279), .B2(n8124), .C1(n7280), .C2(n8060), .A(n7732), 
        .ZN(n7727) );
  OAI222_X1 U6883 ( .A1(n5082), .A2(n7282), .B1(n937), .B2(n5825), .C1(n5485), 
        .C2(n5816), .ZN(n7732) );
  AOI221_X1 U6884 ( .B1(n5833), .B2(DATAIN[56]), .C1(n7283), .C2(OUT2[56]), 
        .A(n7733), .ZN(n7726) );
  OAI22_X1 U6885 ( .A1(n4887), .A2(n5827), .B1(n5421), .B2(n7285), .ZN(n7733)
         );
  NAND4_X1 U6886 ( .A1(n7734), .A2(n7735), .A3(n7736), .A4(n7737), .ZN(n3607)
         );
  AOI221_X1 U6887 ( .B1(n7271), .B2(n5293), .C1(n7272), .C2(n5018), .A(n7738), 
        .ZN(n7737) );
  OAI222_X1 U6888 ( .A1(n1064), .A2(n5820), .B1(n1000), .B2(n5823), .C1(n1128), 
        .C2(n5815), .ZN(n7738) );
  AOI221_X1 U6889 ( .B1(n7274), .B2(n5358), .C1(n7275), .C2(n5147), .A(n7739), 
        .ZN(n7736) );
  OAI222_X1 U6890 ( .A1(n552), .A2(n7277), .B1(n488), .B2(n5824), .C1(n744), 
        .C2(n7278), .ZN(n7739) );
  AOI221_X1 U6891 ( .B1(n7279), .B2(n8123), .C1(n7280), .C2(n8059), .A(n7740), 
        .ZN(n7735) );
  OAI222_X1 U6892 ( .A1(n5083), .A2(n7282), .B1(n936), .B2(n5825), .C1(n5486), 
        .C2(n5816), .ZN(n7740) );
  AOI221_X1 U6893 ( .B1(n5833), .B2(DATAIN[57]), .C1(n7283), .C2(OUT2[57]), 
        .A(n7741), .ZN(n7734) );
  OAI22_X1 U6894 ( .A1(n4888), .A2(n5827), .B1(n5422), .B2(n7285), .ZN(n7741)
         );
  NAND4_X1 U6895 ( .A1(n7742), .A2(n7743), .A3(n7744), .A4(n7745), .ZN(n3606)
         );
  AOI221_X1 U6896 ( .B1(n7271), .B2(n5294), .C1(n7272), .C2(n5019), .A(n7746), 
        .ZN(n7745) );
  OAI222_X1 U6897 ( .A1(n1063), .A2(n5820), .B1(n999), .B2(n5823), .C1(n1127), 
        .C2(n5815), .ZN(n7746) );
  AOI221_X1 U6898 ( .B1(n7274), .B2(n5359), .C1(n7275), .C2(n5148), .A(n7747), 
        .ZN(n7744) );
  OAI222_X1 U6899 ( .A1(n551), .A2(n7277), .B1(n487), .B2(n5824), .C1(n743), 
        .C2(n7278), .ZN(n7747) );
  AOI221_X1 U6900 ( .B1(n7279), .B2(n8122), .C1(n7280), .C2(n8058), .A(n7748), 
        .ZN(n7743) );
  OAI222_X1 U6901 ( .A1(n5084), .A2(n7282), .B1(n935), .B2(n5825), .C1(n5487), 
        .C2(n5816), .ZN(n7748) );
  AOI221_X1 U6902 ( .B1(n5833), .B2(DATAIN[58]), .C1(n7283), .C2(OUT2[58]), 
        .A(n7749), .ZN(n7742) );
  OAI22_X1 U6903 ( .A1(n4889), .A2(n5827), .B1(n5423), .B2(n7285), .ZN(n7749)
         );
  NAND4_X1 U6904 ( .A1(n7750), .A2(n7751), .A3(n7752), .A4(n7753), .ZN(n3605)
         );
  AOI221_X1 U6905 ( .B1(n7271), .B2(n5295), .C1(n7272), .C2(n5020), .A(n7754), 
        .ZN(n7753) );
  OAI222_X1 U6906 ( .A1(n1062), .A2(n5820), .B1(n998), .B2(n5823), .C1(n1126), 
        .C2(n5815), .ZN(n7754) );
  AOI221_X1 U6907 ( .B1(n7274), .B2(n5360), .C1(n7275), .C2(n5149), .A(n7755), 
        .ZN(n7752) );
  OAI222_X1 U6908 ( .A1(n550), .A2(n7277), .B1(n486), .B2(n5824), .C1(n742), 
        .C2(n7278), .ZN(n7755) );
  AOI221_X1 U6909 ( .B1(n7279), .B2(n8121), .C1(n7280), .C2(n8057), .A(n7756), 
        .ZN(n7751) );
  OAI222_X1 U6910 ( .A1(n5085), .A2(n7282), .B1(n934), .B2(n5825), .C1(n5488), 
        .C2(n5816), .ZN(n7756) );
  AOI221_X1 U6911 ( .B1(n5833), .B2(DATAIN[59]), .C1(n7283), .C2(OUT2[59]), 
        .A(n7757), .ZN(n7750) );
  OAI22_X1 U6912 ( .A1(n4890), .A2(n5827), .B1(n5424), .B2(n7285), .ZN(n7757)
         );
  NAND4_X1 U6913 ( .A1(n7758), .A2(n7759), .A3(n7760), .A4(n7761), .ZN(n3604)
         );
  AOI221_X1 U6914 ( .B1(n7271), .B2(n5296), .C1(n7272), .C2(n5021), .A(n7762), 
        .ZN(n7761) );
  OAI222_X1 U6915 ( .A1(n1061), .A2(n5820), .B1(n997), .B2(n5823), .C1(n1125), 
        .C2(n5815), .ZN(n7762) );
  AOI221_X1 U6916 ( .B1(n7274), .B2(n5361), .C1(n7275), .C2(n5150), .A(n7763), 
        .ZN(n7760) );
  OAI222_X1 U6917 ( .A1(n549), .A2(n7277), .B1(n485), .B2(n5824), .C1(n741), 
        .C2(n7278), .ZN(n7763) );
  AOI221_X1 U6918 ( .B1(n7279), .B2(n8120), .C1(n7280), .C2(n8056), .A(n7764), 
        .ZN(n7759) );
  OAI222_X1 U6919 ( .A1(n5086), .A2(n7282), .B1(n933), .B2(n5825), .C1(n5489), 
        .C2(n5816), .ZN(n7764) );
  AOI221_X1 U6920 ( .B1(n5833), .B2(DATAIN[60]), .C1(n7283), .C2(OUT2[60]), 
        .A(n7765), .ZN(n7758) );
  OAI22_X1 U6921 ( .A1(n4891), .A2(n5827), .B1(n5425), .B2(n7285), .ZN(n7765)
         );
  NAND4_X1 U6922 ( .A1(n7766), .A2(n7767), .A3(n7768), .A4(n7769), .ZN(n3603)
         );
  AOI221_X1 U6923 ( .B1(n7271), .B2(n5297), .C1(n7272), .C2(n5022), .A(n7770), 
        .ZN(n7769) );
  OAI222_X1 U6924 ( .A1(n1060), .A2(n5820), .B1(n996), .B2(n5823), .C1(n1124), 
        .C2(n5815), .ZN(n7770) );
  AOI221_X1 U6925 ( .B1(n7274), .B2(n5362), .C1(n7275), .C2(n5151), .A(n7771), 
        .ZN(n7768) );
  OAI222_X1 U6926 ( .A1(n548), .A2(n7277), .B1(n484), .B2(n5824), .C1(n740), 
        .C2(n7278), .ZN(n7771) );
  AOI221_X1 U6927 ( .B1(n7279), .B2(n8119), .C1(n7280), .C2(n8055), .A(n7772), 
        .ZN(n7767) );
  OAI222_X1 U6928 ( .A1(n5087), .A2(n7282), .B1(n932), .B2(n5825), .C1(n5490), 
        .C2(n5816), .ZN(n7772) );
  AOI221_X1 U6929 ( .B1(n5833), .B2(DATAIN[61]), .C1(n7283), .C2(OUT2[61]), 
        .A(n7773), .ZN(n7766) );
  OAI22_X1 U6930 ( .A1(n4892), .A2(n5827), .B1(n5426), .B2(n7285), .ZN(n7773)
         );
  NAND4_X1 U6931 ( .A1(n7774), .A2(n7775), .A3(n7776), .A4(n7777), .ZN(n3602)
         );
  AOI221_X1 U6932 ( .B1(n7271), .B2(n5298), .C1(n7272), .C2(n5023), .A(n7778), 
        .ZN(n7777) );
  OAI222_X1 U6933 ( .A1(n1059), .A2(n5820), .B1(n995), .B2(n5823), .C1(n1123), 
        .C2(n5815), .ZN(n7778) );
  AOI221_X1 U6934 ( .B1(n7274), .B2(n5363), .C1(n7275), .C2(n5152), .A(n7779), 
        .ZN(n7776) );
  OAI222_X1 U6935 ( .A1(n547), .A2(n7277), .B1(n483), .B2(n5824), .C1(n739), 
        .C2(n7278), .ZN(n7779) );
  AOI221_X1 U6936 ( .B1(n7279), .B2(n8118), .C1(n7280), .C2(n8054), .A(n7780), 
        .ZN(n7775) );
  OAI222_X1 U6937 ( .A1(n5088), .A2(n7282), .B1(n931), .B2(n5825), .C1(n5491), 
        .C2(n5816), .ZN(n7780) );
  AOI221_X1 U6938 ( .B1(n5833), .B2(DATAIN[62]), .C1(n7283), .C2(OUT2[62]), 
        .A(n7781), .ZN(n7774) );
  OAI22_X1 U6939 ( .A1(n4893), .A2(n5827), .B1(n5427), .B2(n7285), .ZN(n7781)
         );
  NAND4_X1 U6940 ( .A1(n7782), .A2(n7783), .A3(n7784), .A4(n7785), .ZN(n3601)
         );
  AOI221_X1 U6941 ( .B1(n7271), .B2(n5299), .C1(n7272), .C2(n5024), .A(n7786), 
        .ZN(n7785) );
  OAI222_X1 U6942 ( .A1(n1058), .A2(n5820), .B1(n994), .B2(n5823), .C1(n1122), 
        .C2(n5815), .ZN(n7786) );
  AND3_X1 U6943 ( .A1(N434), .A2(n5852), .A3(N435), .ZN(n7787) );
  AOI221_X1 U6944 ( .B1(n7274), .B2(n5364), .C1(n7275), .C2(n5153), .A(n7795), 
        .ZN(n7784) );
  OAI222_X1 U6945 ( .A1(n546), .A2(n7277), .B1(n482), .B2(n5824), .C1(n738), 
        .C2(n7278), .ZN(n7795) );
  NOR3_X1 U6946 ( .A1(N433), .A2(N434), .A3(n7796), .ZN(n7794) );
  NOR2_X1 U6947 ( .A1(n7789), .A2(n5852), .ZN(n7791) );
  AOI221_X1 U6948 ( .B1(n7279), .B2(n8117), .C1(n7280), .C2(n8053), .A(n7799), 
        .ZN(n7783) );
  OAI222_X1 U6949 ( .A1(n5089), .A2(n7282), .B1(n930), .B2(n5825), .C1(n5492), 
        .C2(n5816), .ZN(n7799) );
  AND2_X1 U6950 ( .A1(n7788), .A2(N435), .ZN(n7790) );
  INV_X1 U6951 ( .A(n7801), .ZN(n7788) );
  AND2_X1 U6952 ( .A1(n7793), .A2(N434), .ZN(n7797) );
  AOI221_X1 U6953 ( .B1(n5833), .B2(DATAIN[63]), .C1(n7283), .C2(OUT2[63]), 
        .A(n7802), .ZN(n7782) );
  OAI22_X1 U6954 ( .A1(n4894), .A2(n5827), .B1(n5428), .B2(n7285), .ZN(n7802)
         );
  NOR3_X1 U6955 ( .A1(n7796), .A2(N434), .A3(n7789), .ZN(n7798) );
  INV_X1 U6956 ( .A(N433), .ZN(n7789) );
  INV_X1 U6957 ( .A(n5852), .ZN(n7796) );
  INV_X1 U6958 ( .A(n5864), .ZN(n7803) );
  INV_X1 U6959 ( .A(N434), .ZN(n7792) );
  NOR2_X1 U6960 ( .A1(n7801), .A2(N435), .ZN(n7793) );
  NAND3_X1 U6961 ( .A1(n7804), .A2(n6455), .A3(n7805), .ZN(n7801) );
  NOR2_X1 U6962 ( .A1(N433), .A2(n5852), .ZN(n7800) );
  NAND4_X1 U6963 ( .A1(n7806), .A2(n7807), .A3(WR), .A4(n7808), .ZN(n7805) );
  NOR3_X1 U6964 ( .A1(n7809), .A2(n7810), .A3(n7811), .ZN(n7808) );
  XOR2_X1 U6965 ( .A(n6598), .B(n5860), .Z(n7811) );
  MUX2_X1 U6966 ( .A(n5858), .B(n7812), .S(n7813), .Z(n6598) );
  INV_X1 U6967 ( .A(n7814), .ZN(n7812) );
  XOR2_X1 U6968 ( .A(n6631), .B(N210), .Z(n7810) );
  MUX2_X1 U6969 ( .A(N562), .B(n7814), .S(n7813), .Z(n6631) );
  XOR2_X1 U6970 ( .A(n6651), .B(n6616), .Z(n7809) );
  INV_X1 U6971 ( .A(n6629), .ZN(n6616) );
  MUX2_X1 U6972 ( .A(n5857), .B(n7815), .S(n7813), .Z(n6629) );
  INV_X1 U6973 ( .A(ADD_WR[0]), .ZN(n7815) );
  INV_X1 U6974 ( .A(n5855), .ZN(n6651) );
  XOR2_X1 U6975 ( .A(n6619), .B(n6644), .Z(n7807) );
  MUX2_X1 U6976 ( .A(N561), .B(n7814), .S(n7813), .Z(n6644) );
  OAI21_X1 U6977 ( .B1(ADD_WR[0]), .B2(ADD_WR[1]), .A(ADD_WR[2]), .ZN(n7814)
         );
  INV_X1 U6978 ( .A(N209), .ZN(n6619) );
  XOR2_X1 U6979 ( .A(N208), .B(n6643), .Z(n7806) );
  INV_X1 U6980 ( .A(n6604), .ZN(n6643) );
  MUX2_X1 U6981 ( .A(N560), .B(n7816), .S(n7813), .Z(n6604) );
  AND2_X1 U6982 ( .A1(ADD_WR[3]), .A2(n7817), .ZN(n7813) );
  OR3_X1 U6983 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n7817) );
  XNOR2_X1 U6984 ( .A(ADD_WR[1]), .B(ADD_WR[0]), .ZN(n7816) );
  NAND2_X1 U6985 ( .A1(n7818), .A2(n6455), .ZN(n7804) );
  INV_X1 U6986 ( .A(RST), .ZN(n6455) );
  NAND2_X1 U6987 ( .A1(RD2), .A2(n6497), .ZN(n7818) );
  INV_X1 U6988 ( .A(n8310), .ZN(\r631/carry[1] ) );
  NAND4_X1 U6989 ( .A1(RET), .A2(n6498), .A3(n6494), .A4(n6491), .ZN(n8310) );
  INV_X1 U6990 ( .A(CALL), .ZN(n6491) );
  NAND4_X1 U6991 ( .A1(n1258), .A2(n1260), .A3(n1259), .A4(n7819), .ZN(n6494)
         );
  NOR2_X1 U6992 ( .A1(n5025), .A2(SWP[4]), .ZN(n7819) );
  AND4_X1 U6993 ( .A1(n7820), .A2(n7821), .A3(n7822), .A4(n7823), .ZN(n6498)
         );
  NOR2_X1 U6994 ( .A1(n7824), .A2(n7825), .ZN(n7823) );
  XOR2_X1 U6995 ( .A(n1303), .B(n1250), .Z(n7825) );
  XOR2_X1 U6996 ( .A(n1318), .B(n1261), .Z(n7824) );
  XOR2_X1 U6997 ( .A(n1259), .B(CWP[2]), .Z(n7822) );
  XOR2_X1 U6998 ( .A(SWP[1]), .B(n1317), .Z(n7821) );
  XOR2_X1 U6999 ( .A(SWP[3]), .B(n1315), .Z(n7820) );
  NOR2_X1 U7000 ( .A1(n7826), .A2(n7827), .ZN(\U3/U202/Z_3 ) );
  INV_X1 U7001 ( .A(\U3/U195/Z_3 ), .ZN(n7826) );
  OAI222_X1 U7002 ( .A1(n7827), .A2(n7828), .B1(n7829), .B2(n7830), .C1(n1328), 
        .C2(n7831), .ZN(\U3/U202/Z_2 ) );
  OAI222_X1 U7003 ( .A1(n7827), .A2(n7832), .B1(n7833), .B2(n7829), .C1(n7831), 
        .C2(n5300), .ZN(\U3/U202/Z_1 ) );
  INV_X1 U7004 ( .A(n7834), .ZN(n7833) );
  OAI21_X1 U7005 ( .B1(n1330), .B2(n7831), .A(n7835), .ZN(\U3/U202/Z_0 ) );
  MUX2_X1 U7006 ( .A(n7829), .B(n7827), .S(ADD_RD2[0]), .Z(n7835) );
  NOR2_X1 U7007 ( .A1(n1303), .A2(n7836), .ZN(\U3/U201/Z_4 ) );
  OAI21_X1 U7008 ( .B1(n1315), .B2(n7836), .A(n7829), .ZN(\U3/U201/Z_3 ) );
  OAI21_X1 U7009 ( .B1(n1316), .B2(n7836), .A(n7829), .ZN(\U3/U201/Z_2 ) );
  NAND2_X1 U7010 ( .A1(n7837), .A2(n6645), .ZN(n7829) );
  NOR2_X1 U7011 ( .A1(n1317), .A2(n7836), .ZN(\U3/U201/Z_1 ) );
  NOR2_X1 U7012 ( .A1(n1318), .A2(n7836), .ZN(\U3/U201/Z_0 ) );
  AND3_X1 U7013 ( .A1(n7827), .A2(n6654), .A3(n1322), .ZN(n7836) );
  NAND2_X1 U7014 ( .A1(n6645), .A2(n7838), .ZN(n7827) );
  INV_X1 U7015 ( .A(n6720), .ZN(n6645) );
  NOR2_X1 U7016 ( .A1(n1303), .A2(n7839), .ZN(\U3/U200/Z_4 ) );
  NOR2_X1 U7017 ( .A1(n1315), .A2(n7839), .ZN(\U3/U200/Z_3 ) );
  INV_X1 U7018 ( .A(n7840), .ZN(\U3/U200/Z_2 ) );
  MUX2_X1 U7019 ( .A(n1316), .B(n6481), .S(n7839), .Z(n7840) );
  MUX2_X1 U7020 ( .A(n7841), .B(n7842), .S(n7843), .Z(n6481) );
  OAI22_X1 U7021 ( .A1(n7844), .A2(n1328), .B1(n7845), .B2(n7846), .ZN(n7843)
         );
  XOR2_X1 U7022 ( .A(n7847), .B(n7848), .Z(n7842) );
  NAND2_X1 U7023 ( .A1(n6479), .A2(n7849), .ZN(n7848) );
  NAND3_X1 U7024 ( .A1(n7849), .A2(n6479), .A3(n7846), .ZN(n7841) );
  MUX2_X1 U7025 ( .A(CWP[1]), .B(n6514), .S(n7839), .Z(\U3/U200/Z_1 ) );
  OAI21_X1 U7026 ( .B1(n7850), .B2(n7851), .A(n7847), .ZN(n6514) );
  NAND2_X1 U7027 ( .A1(n7850), .A2(n7851), .ZN(n7847) );
  XNOR2_X1 U7028 ( .A(n7849), .B(n6479), .ZN(n7850) );
  OAI22_X1 U7029 ( .A1(n7846), .A2(n7852), .B1(n7844), .B2(n5300), .ZN(n7849)
         );
  INV_X1 U7030 ( .A(n7853), .ZN(\U3/U200/Z_0 ) );
  MUX2_X1 U7031 ( .A(n1318), .B(n6479), .S(n7839), .Z(n7853) );
  OAI22_X1 U7032 ( .A1(n7846), .A2(n7854), .B1(n1330), .B2(n7844), .ZN(n6479)
         );
  OAI21_X1 U7033 ( .B1(n6475), .B2(SPILL), .A(n6513), .ZN(n7844) );
  INV_X1 U7034 ( .A(n6476), .ZN(n6513) );
  NOR3_X1 U7035 ( .A1(n1330), .A2(n8309), .A3(n1328), .ZN(n6476) );
  INV_X1 U7036 ( .A(n6654), .ZN(n6475) );
  NAND2_X1 U7037 ( .A1(n1322), .A2(FILL), .ZN(n6654) );
  INV_X1 U7038 ( .A(n7851), .ZN(n7846) );
  NAND2_X1 U7039 ( .A1(n7266), .A2(n6720), .ZN(n7851) );
  NAND2_X1 U7040 ( .A1(WR), .A2(n6497), .ZN(n6720) );
  NAND2_X1 U7041 ( .A1(RD1), .A2(n6497), .ZN(n7266) );
  INV_X1 U7042 ( .A(n6507), .ZN(n6497) );
  NAND2_X1 U7043 ( .A1(EN), .A2(n7831), .ZN(n6507) );
  NOR2_X1 U7044 ( .A1(FILL), .A2(SPILL), .ZN(n7831) );
  NAND2_X1 U7045 ( .A1(n7845), .A2(n7855), .ZN(\U3/U199/Z_2 ) );
  NOR2_X1 U7046 ( .A1(n7839), .A2(n7852), .ZN(\U3/U199/Z_1 ) );
  NOR2_X1 U7047 ( .A1(n7839), .A2(n7854), .ZN(\U3/U199/Z_0 ) );
  INV_X1 U7048 ( .A(n7855), .ZN(n7839) );
  NAND2_X1 U7049 ( .A1(\U3/U199/Z_3 ), .A2(n7856), .ZN(n7855) );
  NAND3_X1 U7050 ( .A1(n7852), .A2(n7845), .A3(n7854), .ZN(n7856) );
  INV_X1 U7051 ( .A(ADD_RD1[0]), .ZN(n7854) );
  INV_X1 U7052 ( .A(ADD_RD1[2]), .ZN(n7845) );
  INV_X1 U7053 ( .A(ADD_RD1[1]), .ZN(n7852) );
  NOR2_X1 U7054 ( .A1(n1303), .A2(n7837), .ZN(\U3/U196/Z_4 ) );
  NOR2_X1 U7055 ( .A1(n1315), .A2(n7837), .ZN(\U3/U196/Z_3 ) );
  INV_X1 U7056 ( .A(n7857), .ZN(\U3/U196/Z_2 ) );
  MUX2_X1 U7057 ( .A(n1316), .B(n7830), .S(n7837), .Z(n7857) );
  NAND2_X1 U7058 ( .A1(ADD_RD2[2]), .A2(n7858), .ZN(n7830) );
  MUX2_X1 U7059 ( .A(CWP[1]), .B(n7834), .S(n7837), .Z(\U3/U196/Z_1 ) );
  OAI21_X1 U7060 ( .B1(n7859), .B2(n7832), .A(n7858), .ZN(n7834) );
  INV_X1 U7061 ( .A(n7860), .ZN(\U3/U196/Z_0 ) );
  MUX2_X1 U7062 ( .A(n1318), .B(ADD_RD2[0]), .S(n7837), .Z(n7860) );
  NAND2_X1 U7063 ( .A1(n7828), .A2(n7838), .ZN(\U3/U195/Z_2 ) );
  INV_X1 U7064 ( .A(ADD_RD2[2]), .ZN(n7828) );
  NOR2_X1 U7065 ( .A1(n7837), .A2(n7832), .ZN(\U3/U195/Z_1 ) );
  NOR2_X1 U7066 ( .A1(n7837), .A2(n7859), .ZN(\U3/U195/Z_0 ) );
  INV_X1 U7067 ( .A(n7838), .ZN(n7837) );
  OAI21_X1 U7068 ( .B1(ADD_RD2[2]), .B2(n7858), .A(\U3/U195/Z_3 ), .ZN(n7838)
         );
  NAND2_X1 U7069 ( .A1(n7859), .A2(n7832), .ZN(n7858) );
  INV_X1 U7070 ( .A(ADD_RD2[1]), .ZN(n7832) );
  INV_X1 U7071 ( .A(ADD_RD2[0]), .ZN(n7859) );
endmodule

