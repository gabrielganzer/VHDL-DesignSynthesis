----------------------------------------------------------------------------------
-- Engineer: GANZER Gabriel
-- Company: Politecnico di Torino
-- File : constants.vhd
-- Descriptions: constants used throughout project
-- Date: 14/04/2020
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package CONSTANTS is 
   constant WIDTH : integer := 32;
   constant STEP : integer := 4;
end package;